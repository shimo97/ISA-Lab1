library verilog;
use verilog.vl_types.all;
entity tb_mul is
end tb_mul;
