library verilog;
use verilog.vl_types.all;
entity tb_fir_LA is
end tb_fir_LA;
