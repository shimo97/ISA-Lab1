LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY DADDA IS
PORT(
Li : IN std_logic_vector(26 downto 0);
Mi : IN std_logic_vector(24 downto 0);
Ki : IN std_logic_vector(27 downto 0);
Ji : IN std_logic_vector(27 downto 0);
Ii : IN std_logic_vector(27 downto 0);
Hi : IN std_logic_vector(27 downto 0);
Gi : IN std_logic_vector(27 downto 0);
Fi : IN std_logic_vector(27 downto 0);
Ei : IN std_logic_vector(27 downto 0);
Di : IN std_logic_vector(27 downto 0);
Ci : IN std_logic_vector(27 downto 0);
Bi : IN std_logic_vector(27 downto 0);
Ai : IN std_logic_vector(27 downto 0);
Y : OUT std_logic_vector(47 downto 0));
END DADDA;

ARCHITECTURE behavior OF DADDA IS

SIGNAL N0_358 : std_logic;
SIGNAL N0_359 : std_logic;
SIGNAL N0_355 : std_logic;
SIGNAL N0_356 : std_logic;
SIGNAL N0_357 : std_logic;
SIGNAL N0_352 : std_logic;
SIGNAL N0_353 : std_logic;
SIGNAL N0_354 : std_logic;
SIGNAL N0_348 : std_logic;
SIGNAL N0_349 : std_logic;
SIGNAL N0_350 : std_logic;
SIGNAL N0_351 : std_logic;
SIGNAL N0_344 : std_logic;
SIGNAL N0_345 : std_logic;
SIGNAL N0_346 : std_logic;
SIGNAL N0_347 : std_logic;
SIGNAL N0_339 : std_logic;
SIGNAL N0_340 : std_logic;
SIGNAL N0_341 : std_logic;
SIGNAL N0_342 : std_logic;
SIGNAL N0_343 : std_logic;
SIGNAL N0_334 : std_logic;
SIGNAL N0_335 : std_logic;
SIGNAL N0_336 : std_logic;
SIGNAL N0_337 : std_logic;
SIGNAL N0_338 : std_logic;
SIGNAL N0_328 : std_logic;
SIGNAL N0_329 : std_logic;
SIGNAL N0_330 : std_logic;
SIGNAL N0_331 : std_logic;
SIGNAL N0_332 : std_logic;
SIGNAL N0_333 : std_logic;
SIGNAL N0_322 : std_logic;
SIGNAL N0_323 : std_logic;
SIGNAL N0_324 : std_logic;
SIGNAL N0_325 : std_logic;
SIGNAL N0_326 : std_logic;
SIGNAL N0_327 : std_logic;
SIGNAL N0_315 : std_logic;
SIGNAL N0_316 : std_logic;
SIGNAL N0_317 : std_logic;
SIGNAL N0_318 : std_logic;
SIGNAL N0_319 : std_logic;
SIGNAL N0_320 : std_logic;
SIGNAL N0_321 : std_logic;
SIGNAL N0_308 : std_logic;
SIGNAL N0_309 : std_logic;
SIGNAL N0_310 : std_logic;
SIGNAL N0_311 : std_logic;
SIGNAL N0_312 : std_logic;
SIGNAL N0_313 : std_logic;
SIGNAL N0_314 : std_logic;
SIGNAL N0_300 : std_logic;
SIGNAL N0_301 : std_logic;
SIGNAL N0_302 : std_logic;
SIGNAL N0_303 : std_logic;
SIGNAL N0_304 : std_logic;
SIGNAL N0_305 : std_logic;
SIGNAL N0_306 : std_logic;
SIGNAL N0_307 : std_logic;
SIGNAL N0_292 : std_logic;
SIGNAL N0_293 : std_logic;
SIGNAL N0_294 : std_logic;
SIGNAL N0_295 : std_logic;
SIGNAL N0_296 : std_logic;
SIGNAL N0_297 : std_logic;
SIGNAL N0_298 : std_logic;
SIGNAL N0_299 : std_logic;
SIGNAL N0_283 : std_logic;
SIGNAL N0_284 : std_logic;
SIGNAL N0_285 : std_logic;
SIGNAL N0_286 : std_logic;
SIGNAL N0_287 : std_logic;
SIGNAL N0_288 : std_logic;
SIGNAL N0_289 : std_logic;
SIGNAL N0_290 : std_logic;
SIGNAL N0_291 : std_logic;
SIGNAL N0_274 : std_logic;
SIGNAL N0_275 : std_logic;
SIGNAL N0_276 : std_logic;
SIGNAL N0_277 : std_logic;
SIGNAL N0_278 : std_logic;
SIGNAL N0_279 : std_logic;
SIGNAL N0_280 : std_logic;
SIGNAL N0_281 : std_logic;
SIGNAL N0_282 : std_logic;
SIGNAL N0_264 : std_logic;
SIGNAL N0_265 : std_logic;
SIGNAL N0_266 : std_logic;
SIGNAL N0_267 : std_logic;
SIGNAL N0_268 : std_logic;
SIGNAL N0_269 : std_logic;
SIGNAL N0_270 : std_logic;
SIGNAL N0_271 : std_logic;
SIGNAL N0_272 : std_logic;
SIGNAL N0_273 : std_logic;
SIGNAL N0_254 : std_logic;
SIGNAL N0_255 : std_logic;
SIGNAL N0_256 : std_logic;
SIGNAL N0_257 : std_logic;
SIGNAL N0_258 : std_logic;
SIGNAL N0_259 : std_logic;
SIGNAL N0_260 : std_logic;
SIGNAL N0_261 : std_logic;
SIGNAL N0_262 : std_logic;
SIGNAL N0_263 : std_logic;
SIGNAL N0_243 : std_logic;
SIGNAL N0_244 : std_logic;
SIGNAL N0_245 : std_logic;
SIGNAL N0_246 : std_logic;
SIGNAL N0_247 : std_logic;
SIGNAL N0_248 : std_logic;
SIGNAL N0_249 : std_logic;
SIGNAL N0_250 : std_logic;
SIGNAL N0_251 : std_logic;
SIGNAL N0_252 : std_logic;
SIGNAL N0_253 : std_logic;
SIGNAL N0_232 : std_logic;
SIGNAL N0_233 : std_logic;
SIGNAL N0_234 : std_logic;
SIGNAL N0_235 : std_logic;
SIGNAL N0_236 : std_logic;
SIGNAL N0_237 : std_logic;
SIGNAL N0_238 : std_logic;
SIGNAL N0_239 : std_logic;
SIGNAL N0_240 : std_logic;
SIGNAL N0_241 : std_logic;
SIGNAL N0_242 : std_logic;
SIGNAL N0_220 : std_logic;
SIGNAL N0_221 : std_logic;
SIGNAL N0_222 : std_logic;
SIGNAL N0_223 : std_logic;
SIGNAL N0_224 : std_logic;
SIGNAL N0_225 : std_logic;
SIGNAL N0_226 : std_logic;
SIGNAL N0_227 : std_logic;
SIGNAL N0_228 : std_logic;
SIGNAL N0_229 : std_logic;
SIGNAL N0_230 : std_logic;
SIGNAL N0_231 : std_logic;
SIGNAL N0_207 : std_logic;
SIGNAL N0_208 : std_logic;
SIGNAL N0_209 : std_logic;
SIGNAL N0_210 : std_logic;
SIGNAL N0_211 : std_logic;
SIGNAL N0_212 : std_logic;
SIGNAL N0_213 : std_logic;
SIGNAL N0_214 : std_logic;
SIGNAL N0_215 : std_logic;
SIGNAL N0_216 : std_logic;
SIGNAL N0_217 : std_logic;
SIGNAL N0_218 : std_logic;
SIGNAL N0_219 : std_logic;
SIGNAL N0_194 : std_logic;
SIGNAL N0_195 : std_logic;
SIGNAL N0_196 : std_logic;
SIGNAL N0_197 : std_logic;
SIGNAL N0_198 : std_logic;
SIGNAL N0_199 : std_logic;
SIGNAL N0_200 : std_logic;
SIGNAL N0_201 : std_logic;
SIGNAL N0_202 : std_logic;
SIGNAL N0_203 : std_logic;
SIGNAL N0_204 : std_logic;
SIGNAL N0_205 : std_logic;
SIGNAL N0_206 : std_logic;
SIGNAL N0_181 : std_logic;
SIGNAL N0_182 : std_logic;
SIGNAL N0_183 : std_logic;
SIGNAL N0_184 : std_logic;
SIGNAL N0_185 : std_logic;
SIGNAL N0_186 : std_logic;
SIGNAL N0_187 : std_logic;
SIGNAL N0_188 : std_logic;
SIGNAL N0_189 : std_logic;
SIGNAL N0_190 : std_logic;
SIGNAL N0_191 : std_logic;
SIGNAL N0_192 : std_logic;
SIGNAL N0_193 : std_logic;
SIGNAL N0_168 : std_logic;
SIGNAL N0_169 : std_logic;
SIGNAL N0_170 : std_logic;
SIGNAL N0_171 : std_logic;
SIGNAL N0_172 : std_logic;
SIGNAL N0_173 : std_logic;
SIGNAL N0_174 : std_logic;
SIGNAL N0_175 : std_logic;
SIGNAL N0_176 : std_logic;
SIGNAL N0_177 : std_logic;
SIGNAL N0_178 : std_logic;
SIGNAL N0_179 : std_logic;
SIGNAL N0_180 : std_logic;
SIGNAL N0_156 : std_logic;
SIGNAL N0_157 : std_logic;
SIGNAL N0_158 : std_logic;
SIGNAL N0_159 : std_logic;
SIGNAL N0_160 : std_logic;
SIGNAL N0_161 : std_logic;
SIGNAL N0_162 : std_logic;
SIGNAL N0_163 : std_logic;
SIGNAL N0_164 : std_logic;
SIGNAL N0_165 : std_logic;
SIGNAL N0_166 : std_logic;
SIGNAL N0_167 : std_logic;
SIGNAL N0_143 : std_logic;
SIGNAL N0_144 : std_logic;
SIGNAL N0_145 : std_logic;
SIGNAL N0_146 : std_logic;
SIGNAL N0_147 : std_logic;
SIGNAL N0_148 : std_logic;
SIGNAL N0_149 : std_logic;
SIGNAL N0_150 : std_logic;
SIGNAL N0_151 : std_logic;
SIGNAL N0_152 : std_logic;
SIGNAL N0_153 : std_logic;
SIGNAL N0_154 : std_logic;
SIGNAL N0_155 : std_logic;
SIGNAL N0_132 : std_logic;
SIGNAL N0_133 : std_logic;
SIGNAL N0_134 : std_logic;
SIGNAL N0_135 : std_logic;
SIGNAL N0_136 : std_logic;
SIGNAL N0_137 : std_logic;
SIGNAL N0_138 : std_logic;
SIGNAL N0_139 : std_logic;
SIGNAL N0_140 : std_logic;
SIGNAL N0_141 : std_logic;
SIGNAL N0_142 : std_logic;
SIGNAL N0_120 : std_logic;
SIGNAL N0_121 : std_logic;
SIGNAL N0_122 : std_logic;
SIGNAL N0_123 : std_logic;
SIGNAL N0_124 : std_logic;
SIGNAL N0_125 : std_logic;
SIGNAL N0_126 : std_logic;
SIGNAL N0_127 : std_logic;
SIGNAL N0_128 : std_logic;
SIGNAL N0_129 : std_logic;
SIGNAL N0_130 : std_logic;
SIGNAL N0_131 : std_logic;
SIGNAL N0_110 : std_logic;
SIGNAL N0_111 : std_logic;
SIGNAL N0_112 : std_logic;
SIGNAL N0_113 : std_logic;
SIGNAL N0_114 : std_logic;
SIGNAL N0_115 : std_logic;
SIGNAL N0_116 : std_logic;
SIGNAL N0_117 : std_logic;
SIGNAL N0_118 : std_logic;
SIGNAL N0_119 : std_logic;
SIGNAL N0_99 : std_logic;
SIGNAL N0_100 : std_logic;
SIGNAL N0_101 : std_logic;
SIGNAL N0_102 : std_logic;
SIGNAL N0_103 : std_logic;
SIGNAL N0_104 : std_logic;
SIGNAL N0_105 : std_logic;
SIGNAL N0_106 : std_logic;
SIGNAL N0_107 : std_logic;
SIGNAL N0_108 : std_logic;
SIGNAL N0_109 : std_logic;
SIGNAL N0_90 : std_logic;
SIGNAL N0_91 : std_logic;
SIGNAL N0_92 : std_logic;
SIGNAL N0_93 : std_logic;
SIGNAL N0_94 : std_logic;
SIGNAL N0_95 : std_logic;
SIGNAL N0_96 : std_logic;
SIGNAL N0_97 : std_logic;
SIGNAL N0_98 : std_logic;
SIGNAL N0_80 : std_logic;
SIGNAL N0_81 : std_logic;
SIGNAL N0_82 : std_logic;
SIGNAL N0_83 : std_logic;
SIGNAL N0_84 : std_logic;
SIGNAL N0_85 : std_logic;
SIGNAL N0_86 : std_logic;
SIGNAL N0_87 : std_logic;
SIGNAL N0_88 : std_logic;
SIGNAL N0_89 : std_logic;
SIGNAL N0_72 : std_logic;
SIGNAL N0_73 : std_logic;
SIGNAL N0_74 : std_logic;
SIGNAL N0_75 : std_logic;
SIGNAL N0_76 : std_logic;
SIGNAL N0_77 : std_logic;
SIGNAL N0_78 : std_logic;
SIGNAL N0_79 : std_logic;
SIGNAL N0_63 : std_logic;
SIGNAL N0_64 : std_logic;
SIGNAL N0_65 : std_logic;
SIGNAL N0_66 : std_logic;
SIGNAL N0_67 : std_logic;
SIGNAL N0_68 : std_logic;
SIGNAL N0_69 : std_logic;
SIGNAL N0_70 : std_logic;
SIGNAL N0_71 : std_logic;
SIGNAL N0_56 : std_logic;
SIGNAL N0_57 : std_logic;
SIGNAL N0_58 : std_logic;
SIGNAL N0_59 : std_logic;
SIGNAL N0_60 : std_logic;
SIGNAL N0_61 : std_logic;
SIGNAL N0_62 : std_logic;
SIGNAL N0_48 : std_logic;
SIGNAL N0_49 : std_logic;
SIGNAL N0_50 : std_logic;
SIGNAL N0_51 : std_logic;
SIGNAL N0_52 : std_logic;
SIGNAL N0_53 : std_logic;
SIGNAL N0_54 : std_logic;
SIGNAL N0_55 : std_logic;
SIGNAL N0_42 : std_logic;
SIGNAL N0_43 : std_logic;
SIGNAL N0_44 : std_logic;
SIGNAL N0_45 : std_logic;
SIGNAL N0_46 : std_logic;
SIGNAL N0_47 : std_logic;
SIGNAL N0_35 : std_logic;
SIGNAL N0_36 : std_logic;
SIGNAL N0_37 : std_logic;
SIGNAL N0_38 : std_logic;
SIGNAL N0_39 : std_logic;
SIGNAL N0_40 : std_logic;
SIGNAL N0_41 : std_logic;
SIGNAL N0_30 : std_logic;
SIGNAL N0_31 : std_logic;
SIGNAL N0_32 : std_logic;
SIGNAL N0_33 : std_logic;
SIGNAL N0_34 : std_logic;
SIGNAL N0_24 : std_logic;
SIGNAL N0_25 : std_logic;
SIGNAL N0_26 : std_logic;
SIGNAL N0_27 : std_logic;
SIGNAL N0_28 : std_logic;
SIGNAL N0_29 : std_logic;
SIGNAL N0_20 : std_logic;
SIGNAL N0_21 : std_logic;
SIGNAL N0_22 : std_logic;
SIGNAL N0_23 : std_logic;
SIGNAL N0_15 : std_logic;
SIGNAL N0_16 : std_logic;
SIGNAL N0_17 : std_logic;
SIGNAL N0_18 : std_logic;
SIGNAL N0_19 : std_logic;
SIGNAL N0_12 : std_logic;
SIGNAL N0_13 : std_logic;
SIGNAL N0_14 : std_logic;
SIGNAL N0_8 : std_logic;
SIGNAL N0_9 : std_logic;
SIGNAL N0_10 : std_logic;
SIGNAL N0_11 : std_logic;
SIGNAL N0_6 : std_logic;
SIGNAL N0_7 : std_logic;
SIGNAL N0_3 : std_logic;
SIGNAL N0_4 : std_logic;
SIGNAL N0_5 : std_logic;
SIGNAL N0_2 : std_logic;
SIGNAL N0_0 : std_logic;
SIGNAL N0_1 : std_logic;
SIGNAL N1_0 : std_logic;
SIGNAL N1_1 : std_logic;
SIGNAL N1_2 : std_logic;
SIGNAL N1_3 : std_logic;
SIGNAL N1_4 : std_logic;
SIGNAL N1_5 : std_logic;
SIGNAL N1_6 : std_logic;
SIGNAL N1_7 : std_logic;
SIGNAL N1_8 : std_logic;
SIGNAL N1_9 : std_logic;
SIGNAL N1_10 : std_logic;
SIGNAL N1_11 : std_logic;
SIGNAL N1_12 : std_logic;
SIGNAL N1_13 : std_logic;
SIGNAL N1_14 : std_logic;
SIGNAL N1_15 : std_logic;
SIGNAL N1_16 : std_logic;
SIGNAL N1_17 : std_logic;
SIGNAL N1_18 : std_logic;
SIGNAL N1_19 : std_logic;
SIGNAL N1_20 : std_logic;
SIGNAL N1_21 : std_logic;
SIGNAL N1_22 : std_logic;
SIGNAL N1_23 : std_logic;
SIGNAL N1_24 : std_logic;
SIGNAL N1_25 : std_logic;
SIGNAL N1_26 : std_logic;
SIGNAL N1_27 : std_logic;
SIGNAL N1_28 : std_logic;
SIGNAL N1_29 : std_logic;
SIGNAL N1_30 : std_logic;
SIGNAL N1_31 : std_logic;
SIGNAL N1_32 : std_logic;
SIGNAL N1_33 : std_logic;
SIGNAL N1_34 : std_logic;
SIGNAL N1_35 : std_logic;
SIGNAL N1_36 : std_logic;
SIGNAL N1_37 : std_logic;
SIGNAL N1_38 : std_logic;
SIGNAL N1_39 : std_logic;
SIGNAL N1_40 : std_logic;
SIGNAL N1_41 : std_logic;
SIGNAL N1_42 : std_logic;
SIGNAL N1_43 : std_logic;
SIGNAL N1_44 : std_logic;
SIGNAL N1_45 : std_logic;
SIGNAL N1_46 : std_logic;
SIGNAL N1_47 : std_logic;
SIGNAL N1_48 : std_logic;
SIGNAL N1_49 : std_logic;
SIGNAL N1_50 : std_logic;
SIGNAL N1_51 : std_logic;
SIGNAL N1_52 : std_logic;
SIGNAL N1_53 : std_logic;
SIGNAL N1_54 : std_logic;
SIGNAL N1_55 : std_logic;
SIGNAL N1_56 : std_logic;
SIGNAL N1_57 : std_logic;
SIGNAL N1_58 : std_logic;
SIGNAL N1_59 : std_logic;
SIGNAL N1_60 : std_logic;
SIGNAL N1_61 : std_logic;
SIGNAL N1_62 : std_logic;
SIGNAL N1_63 : std_logic;
SIGNAL N1_64 : std_logic;
SIGNAL N1_65 : std_logic;
SIGNAL N1_66 : std_logic;
SIGNAL N1_67 : std_logic;
SIGNAL N1_68 : std_logic;
SIGNAL N1_69 : std_logic;
SIGNAL N1_70 : std_logic;
SIGNAL N1_71 : std_logic;
SIGNAL N1_72 : std_logic;
SIGNAL N1_73 : std_logic;
SIGNAL N1_74 : std_logic;
SIGNAL N1_75 : std_logic;
SIGNAL N1_76 : std_logic;
SIGNAL N1_77 : std_logic;
SIGNAL N1_78 : std_logic;
SIGNAL N1_79 : std_logic;
SIGNAL H1_0 : std_logic;
SIGNAL C1_0 : std_logic;
SIGNAL N1_80 : std_logic;
SIGNAL N1_81 : std_logic;
SIGNAL N1_82 : std_logic;
SIGNAL N1_83 : std_logic;
SIGNAL N1_84 : std_logic;
SIGNAL N1_85 : std_logic;
SIGNAL N1_86 : std_logic;
SIGNAL N1_87 : std_logic;
SIGNAL H1_1 : std_logic;
SIGNAL C1_1 : std_logic;
SIGNAL N1_88 : std_logic;
SIGNAL N1_89 : std_logic;
SIGNAL N1_90 : std_logic;
SIGNAL N1_91 : std_logic;
SIGNAL N1_92 : std_logic;
SIGNAL N1_93 : std_logic;
SIGNAL N1_94 : std_logic;
SIGNAL F1_0 : std_logic;
SIGNAL C1_2 : std_logic;
SIGNAL H1_2 : std_logic;
SIGNAL C1_3 : std_logic;
SIGNAL N1_95 : std_logic;
SIGNAL N1_96 : std_logic;
SIGNAL N1_97 : std_logic;
SIGNAL N1_98 : std_logic;
SIGNAL N1_99 : std_logic;
SIGNAL N1_100 : std_logic;
SIGNAL F1_1 : std_logic;
SIGNAL C1_4 : std_logic;
SIGNAL H1_3 : std_logic;
SIGNAL C1_5 : std_logic;
SIGNAL N1_101 : std_logic;
SIGNAL N1_102 : std_logic;
SIGNAL N1_103 : std_logic;
SIGNAL N1_104 : std_logic;
SIGNAL N1_105 : std_logic;
SIGNAL F1_2 : std_logic;
SIGNAL C1_6 : std_logic;
SIGNAL F1_3 : std_logic;
SIGNAL C1_7 : std_logic;
SIGNAL H1_4 : std_logic;
SIGNAL C1_8 : std_logic;
SIGNAL N1_106 : std_logic;
SIGNAL N1_107 : std_logic;
SIGNAL N1_108 : std_logic;
SIGNAL N1_109 : std_logic;
SIGNAL F1_4 : std_logic;
SIGNAL C1_9 : std_logic;
SIGNAL F1_5 : std_logic;
SIGNAL C1_10 : std_logic;
SIGNAL H1_5 : std_logic;
SIGNAL C1_11 : std_logic;
SIGNAL N1_110 : std_logic;
SIGNAL N1_111 : std_logic;
SIGNAL N1_112 : std_logic;
SIGNAL F1_6 : std_logic;
SIGNAL C1_12 : std_logic;
SIGNAL F1_7 : std_logic;
SIGNAL C1_13 : std_logic;
SIGNAL F1_8 : std_logic;
SIGNAL C1_14 : std_logic;
SIGNAL H1_6 : std_logic;
SIGNAL C1_15 : std_logic;
SIGNAL N1_113 : std_logic;
SIGNAL N1_114 : std_logic;
SIGNAL F1_9 : std_logic;
SIGNAL C1_16 : std_logic;
SIGNAL F1_10 : std_logic;
SIGNAL C1_17 : std_logic;
SIGNAL F1_11 : std_logic;
SIGNAL C1_18 : std_logic;
SIGNAL H1_7 : std_logic;
SIGNAL C1_19 : std_logic;
SIGNAL N1_115 : std_logic;
SIGNAL F1_12 : std_logic;
SIGNAL C1_20 : std_logic;
SIGNAL F1_13 : std_logic;
SIGNAL C1_21 : std_logic;
SIGNAL F1_14 : std_logic;
SIGNAL C1_22 : std_logic;
SIGNAL F1_15 : std_logic;
SIGNAL C1_23 : std_logic;
SIGNAL N1_116 : std_logic;
SIGNAL F1_16 : std_logic;
SIGNAL C1_24 : std_logic;
SIGNAL F1_17 : std_logic;
SIGNAL C1_25 : std_logic;
SIGNAL F1_18 : std_logic;
SIGNAL C1_26 : std_logic;
SIGNAL F1_19 : std_logic;
SIGNAL C1_27 : std_logic;
SIGNAL N1_117 : std_logic;
SIGNAL F1_20 : std_logic;
SIGNAL C1_28 : std_logic;
SIGNAL F1_21 : std_logic;
SIGNAL C1_29 : std_logic;
SIGNAL F1_22 : std_logic;
SIGNAL C1_30 : std_logic;
SIGNAL F1_23 : std_logic;
SIGNAL C1_31 : std_logic;
SIGNAL N1_118 : std_logic;
SIGNAL F1_24 : std_logic;
SIGNAL C1_32 : std_logic;
SIGNAL F1_25 : std_logic;
SIGNAL C1_33 : std_logic;
SIGNAL F1_26 : std_logic;
SIGNAL C1_34 : std_logic;
SIGNAL F1_27 : std_logic;
SIGNAL C1_35 : std_logic;
SIGNAL N1_119 : std_logic;
SIGNAL F1_28 : std_logic;
SIGNAL C1_36 : std_logic;
SIGNAL F1_29 : std_logic;
SIGNAL C1_37 : std_logic;
SIGNAL F1_30 : std_logic;
SIGNAL C1_38 : std_logic;
SIGNAL H1_8 : std_logic;
SIGNAL C1_39 : std_logic;
SIGNAL N1_120 : std_logic;
SIGNAL F1_31 : std_logic;
SIGNAL C1_40 : std_logic;
SIGNAL F1_32 : std_logic;
SIGNAL C1_41 : std_logic;
SIGNAL F1_33 : std_logic;
SIGNAL C1_42 : std_logic;
SIGNAL N1_121 : std_logic;
SIGNAL N1_122 : std_logic;
SIGNAL F1_34 : std_logic;
SIGNAL C1_43 : std_logic;
SIGNAL F1_35 : std_logic;
SIGNAL C1_44 : std_logic;
SIGNAL H1_9 : std_logic;
SIGNAL C1_45 : std_logic;
SIGNAL N1_123 : std_logic;
SIGNAL N1_124 : std_logic;
SIGNAL N1_125 : std_logic;
SIGNAL F1_36 : std_logic;
SIGNAL C1_46 : std_logic;
SIGNAL F1_37 : std_logic;
SIGNAL C1_47 : std_logic;
SIGNAL N1_126 : std_logic;
SIGNAL N1_127 : std_logic;
SIGNAL N1_128 : std_logic;
SIGNAL N1_129 : std_logic;
SIGNAL F1_38 : std_logic;
SIGNAL C1_48 : std_logic;
SIGNAL H1_10 : std_logic;
SIGNAL C1_49 : std_logic;
SIGNAL N1_130 : std_logic;
SIGNAL N1_131 : std_logic;
SIGNAL N1_132 : std_logic;
SIGNAL N1_133 : std_logic;
SIGNAL N1_134 : std_logic;
SIGNAL F1_39 : std_logic;
SIGNAL C1_50 : std_logic;
SIGNAL N1_135 : std_logic;
SIGNAL N1_136 : std_logic;
SIGNAL N1_137 : std_logic;
SIGNAL N1_138 : std_logic;
SIGNAL N1_139 : std_logic;
SIGNAL N1_140 : std_logic;
SIGNAL H1_11 : std_logic;
SIGNAL C1_51 : std_logic;
SIGNAL N1_141 : std_logic;
SIGNAL N1_142 : std_logic;
SIGNAL N1_143 : std_logic;
SIGNAL N1_144 : std_logic;
SIGNAL N1_145 : std_logic;
SIGNAL N1_146 : std_logic;
SIGNAL N1_147 : std_logic;
SIGNAL N1_148 : std_logic;
SIGNAL N1_149 : std_logic;
SIGNAL N1_150 : std_logic;
SIGNAL N1_151 : std_logic;
SIGNAL N1_152 : std_logic;
SIGNAL N1_153 : std_logic;
SIGNAL N1_154 : std_logic;
SIGNAL N1_155 : std_logic;
SIGNAL N1_156 : std_logic;
SIGNAL N1_157 : std_logic;
SIGNAL N1_158 : std_logic;
SIGNAL N1_159 : std_logic;
SIGNAL N1_160 : std_logic;
SIGNAL N1_161 : std_logic;
SIGNAL N1_162 : std_logic;
SIGNAL N1_163 : std_logic;
SIGNAL N1_164 : std_logic;
SIGNAL N1_165 : std_logic;
SIGNAL N1_166 : std_logic;
SIGNAL N1_167 : std_logic;
SIGNAL N1_168 : std_logic;
SIGNAL N1_169 : std_logic;
SIGNAL N1_170 : std_logic;
SIGNAL N1_171 : std_logic;
SIGNAL N1_172 : std_logic;
SIGNAL N1_173 : std_logic;
SIGNAL N1_174 : std_logic;
SIGNAL N1_175 : std_logic;
SIGNAL N1_176 : std_logic;
SIGNAL N1_177 : std_logic;
SIGNAL N1_178 : std_logic;
SIGNAL N1_179 : std_logic;
SIGNAL N1_180 : std_logic;
SIGNAL N1_181 : std_logic;
SIGNAL N1_182 : std_logic;
SIGNAL N1_183 : std_logic;
SIGNAL N1_184 : std_logic;
SIGNAL N1_185 : std_logic;
SIGNAL N1_186 : std_logic;
SIGNAL N1_187 : std_logic;
SIGNAL N1_188 : std_logic;
SIGNAL N1_189 : std_logic;
SIGNAL N1_190 : std_logic;
SIGNAL N1_191 : std_logic;
SIGNAL N1_192 : std_logic;
SIGNAL N1_193 : std_logic;
SIGNAL N1_194 : std_logic;
SIGNAL N1_195 : std_logic;
SIGNAL N1_196 : std_logic;
SIGNAL N1_197 : std_logic;
SIGNAL N1_198 : std_logic;
SIGNAL N1_199 : std_logic;
SIGNAL N1_200 : std_logic;
SIGNAL N1_201 : std_logic;
SIGNAL N1_202 : std_logic;
SIGNAL N1_203 : std_logic;
SIGNAL N1_204 : std_logic;
SIGNAL N1_205 : std_logic;
SIGNAL N1_206 : std_logic;
SIGNAL N1_207 : std_logic;
SIGNAL N1_208 : std_logic;
SIGNAL N1_209 : std_logic;
SIGNAL N1_210 : std_logic;
SIGNAL N1_211 : std_logic;
SIGNAL N1_212 : std_logic;
SIGNAL N1_213 : std_logic;
SIGNAL N1_214 : std_logic;
SIGNAL N1_215 : std_logic;
SIGNAL N2_0 : std_logic;
SIGNAL N2_1 : std_logic;
SIGNAL N2_2 : std_logic;
SIGNAL N2_3 : std_logic;
SIGNAL N2_4 : std_logic;
SIGNAL N2_5 : std_logic;
SIGNAL N2_6 : std_logic;
SIGNAL N2_7 : std_logic;
SIGNAL N2_8 : std_logic;
SIGNAL N2_9 : std_logic;
SIGNAL N2_10 : std_logic;
SIGNAL N2_11 : std_logic;
SIGNAL N2_12 : std_logic;
SIGNAL N2_13 : std_logic;
SIGNAL N2_14 : std_logic;
SIGNAL N2_15 : std_logic;
SIGNAL N2_16 : std_logic;
SIGNAL N2_17 : std_logic;
SIGNAL N2_18 : std_logic;
SIGNAL N2_19 : std_logic;
SIGNAL N2_20 : std_logic;
SIGNAL N2_21 : std_logic;
SIGNAL N2_22 : std_logic;
SIGNAL N2_23 : std_logic;
SIGNAL N2_24 : std_logic;
SIGNAL N2_25 : std_logic;
SIGNAL N2_26 : std_logic;
SIGNAL N2_27 : std_logic;
SIGNAL N2_28 : std_logic;
SIGNAL N2_29 : std_logic;
SIGNAL N2_30 : std_logic;
SIGNAL N2_31 : std_logic;
SIGNAL N2_32 : std_logic;
SIGNAL N2_33 : std_logic;
SIGNAL N2_34 : std_logic;
SIGNAL H2_0 : std_logic;
SIGNAL C2_0 : std_logic;
SIGNAL N2_35 : std_logic;
SIGNAL N2_36 : std_logic;
SIGNAL N2_37 : std_logic;
SIGNAL N2_38 : std_logic;
SIGNAL N2_39 : std_logic;
SIGNAL H2_1 : std_logic;
SIGNAL C2_1 : std_logic;
SIGNAL N2_40 : std_logic;
SIGNAL N2_41 : std_logic;
SIGNAL N2_42 : std_logic;
SIGNAL N2_43 : std_logic;
SIGNAL F2_0 : std_logic;
SIGNAL C2_2 : std_logic;
SIGNAL H2_2 : std_logic;
SIGNAL C2_3 : std_logic;
SIGNAL N2_44 : std_logic;
SIGNAL N2_45 : std_logic;
SIGNAL N2_46 : std_logic;
SIGNAL F2_1 : std_logic;
SIGNAL C2_4 : std_logic;
SIGNAL H2_3 : std_logic;
SIGNAL C2_5 : std_logic;
SIGNAL N2_47 : std_logic;
SIGNAL N2_48 : std_logic;
SIGNAL F2_2 : std_logic;
SIGNAL C2_6 : std_logic;
SIGNAL F2_3 : std_logic;
SIGNAL C2_7 : std_logic;
SIGNAL H2_4 : std_logic;
SIGNAL C2_8 : std_logic;
SIGNAL N2_49 : std_logic;
SIGNAL F2_4 : std_logic;
SIGNAL C2_9 : std_logic;
SIGNAL F2_5 : std_logic;
SIGNAL C2_10 : std_logic;
SIGNAL H2_5 : std_logic;
SIGNAL C2_11 : std_logic;
SIGNAL F2_6 : std_logic;
SIGNAL C2_12 : std_logic;
SIGNAL F2_7 : std_logic;
SIGNAL C2_13 : std_logic;
SIGNAL F2_8 : std_logic;
SIGNAL C2_14 : std_logic;
SIGNAL F2_9 : std_logic;
SIGNAL C2_15 : std_logic;
SIGNAL F2_10 : std_logic;
SIGNAL C2_16 : std_logic;
SIGNAL F2_11 : std_logic;
SIGNAL C2_17 : std_logic;
SIGNAL F2_12 : std_logic;
SIGNAL C2_18 : std_logic;
SIGNAL F2_13 : std_logic;
SIGNAL C2_19 : std_logic;
SIGNAL F2_14 : std_logic;
SIGNAL C2_20 : std_logic;
SIGNAL F2_15 : std_logic;
SIGNAL C2_21 : std_logic;
SIGNAL F2_16 : std_logic;
SIGNAL C2_22 : std_logic;
SIGNAL F2_17 : std_logic;
SIGNAL C2_23 : std_logic;
SIGNAL F2_18 : std_logic;
SIGNAL C2_24 : std_logic;
SIGNAL F2_19 : std_logic;
SIGNAL C2_25 : std_logic;
SIGNAL F2_20 : std_logic;
SIGNAL C2_26 : std_logic;
SIGNAL F2_21 : std_logic;
SIGNAL C2_27 : std_logic;
SIGNAL F2_22 : std_logic;
SIGNAL C2_28 : std_logic;
SIGNAL F2_23 : std_logic;
SIGNAL C2_29 : std_logic;
SIGNAL F2_24 : std_logic;
SIGNAL C2_30 : std_logic;
SIGNAL F2_25 : std_logic;
SIGNAL C2_31 : std_logic;
SIGNAL F2_26 : std_logic;
SIGNAL C2_32 : std_logic;
SIGNAL F2_27 : std_logic;
SIGNAL C2_33 : std_logic;
SIGNAL F2_28 : std_logic;
SIGNAL C2_34 : std_logic;
SIGNAL F2_29 : std_logic;
SIGNAL C2_35 : std_logic;
SIGNAL F2_30 : std_logic;
SIGNAL C2_36 : std_logic;
SIGNAL F2_31 : std_logic;
SIGNAL C2_37 : std_logic;
SIGNAL F2_32 : std_logic;
SIGNAL C2_38 : std_logic;
SIGNAL F2_33 : std_logic;
SIGNAL C2_39 : std_logic;
SIGNAL F2_34 : std_logic;
SIGNAL C2_40 : std_logic;
SIGNAL F2_35 : std_logic;
SIGNAL C2_41 : std_logic;
SIGNAL F2_36 : std_logic;
SIGNAL C2_42 : std_logic;
SIGNAL F2_37 : std_logic;
SIGNAL C2_43 : std_logic;
SIGNAL F2_38 : std_logic;
SIGNAL C2_44 : std_logic;
SIGNAL F2_39 : std_logic;
SIGNAL C2_45 : std_logic;
SIGNAL F2_40 : std_logic;
SIGNAL C2_46 : std_logic;
SIGNAL F2_41 : std_logic;
SIGNAL C2_47 : std_logic;
SIGNAL F2_42 : std_logic;
SIGNAL C2_48 : std_logic;
SIGNAL F2_43 : std_logic;
SIGNAL C2_49 : std_logic;
SIGNAL F2_44 : std_logic;
SIGNAL C2_50 : std_logic;
SIGNAL F2_45 : std_logic;
SIGNAL C2_51 : std_logic;
SIGNAL F2_46 : std_logic;
SIGNAL C2_52 : std_logic;
SIGNAL F2_47 : std_logic;
SIGNAL C2_53 : std_logic;
SIGNAL F2_48 : std_logic;
SIGNAL C2_54 : std_logic;
SIGNAL F2_49 : std_logic;
SIGNAL C2_55 : std_logic;
SIGNAL F2_50 : std_logic;
SIGNAL C2_56 : std_logic;
SIGNAL F2_51 : std_logic;
SIGNAL C2_57 : std_logic;
SIGNAL F2_52 : std_logic;
SIGNAL C2_58 : std_logic;
SIGNAL F2_53 : std_logic;
SIGNAL C2_59 : std_logic;
SIGNAL F2_54 : std_logic;
SIGNAL C2_60 : std_logic;
SIGNAL F2_55 : std_logic;
SIGNAL C2_61 : std_logic;
SIGNAL F2_56 : std_logic;
SIGNAL C2_62 : std_logic;
SIGNAL F2_57 : std_logic;
SIGNAL C2_63 : std_logic;
SIGNAL F2_58 : std_logic;
SIGNAL C2_64 : std_logic;
SIGNAL F2_59 : std_logic;
SIGNAL C2_65 : std_logic;
SIGNAL F2_60 : std_logic;
SIGNAL C2_66 : std_logic;
SIGNAL F2_61 : std_logic;
SIGNAL C2_67 : std_logic;
SIGNAL F2_62 : std_logic;
SIGNAL C2_68 : std_logic;
SIGNAL F2_63 : std_logic;
SIGNAL C2_69 : std_logic;
SIGNAL F2_64 : std_logic;
SIGNAL C2_70 : std_logic;
SIGNAL F2_65 : std_logic;
SIGNAL C2_71 : std_logic;
SIGNAL F2_66 : std_logic;
SIGNAL C2_72 : std_logic;
SIGNAL F2_67 : std_logic;
SIGNAL C2_73 : std_logic;
SIGNAL H2_6 : std_logic;
SIGNAL C2_74 : std_logic;
SIGNAL F2_68 : std_logic;
SIGNAL C2_75 : std_logic;
SIGNAL F2_69 : std_logic;
SIGNAL C2_76 : std_logic;
SIGNAL N2_50 : std_logic;
SIGNAL F2_70 : std_logic;
SIGNAL C2_77 : std_logic;
SIGNAL H2_7 : std_logic;
SIGNAL C2_78 : std_logic;
SIGNAL N2_51 : std_logic;
SIGNAL N2_52 : std_logic;
SIGNAL F2_71 : std_logic;
SIGNAL C2_79 : std_logic;
SIGNAL N2_53 : std_logic;
SIGNAL N2_54 : std_logic;
SIGNAL N2_55 : std_logic;
SIGNAL H2_8 : std_logic;
SIGNAL C2_80 : std_logic;
SIGNAL N2_56 : std_logic;
SIGNAL N2_57 : std_logic;
SIGNAL N2_58 : std_logic;
SIGNAL N2_59 : std_logic;
SIGNAL N2_60 : std_logic;
SIGNAL N2_61 : std_logic;
SIGNAL N2_62 : std_logic;
SIGNAL N2_63 : std_logic;
SIGNAL N2_64 : std_logic;
SIGNAL N2_65 : std_logic;
SIGNAL N2_66 : std_logic;
SIGNAL N2_67 : std_logic;
SIGNAL N2_68 : std_logic;
SIGNAL N2_69 : std_logic;
SIGNAL N2_70 : std_logic;
SIGNAL N2_71 : std_logic;
SIGNAL N2_72 : std_logic;
SIGNAL N2_73 : std_logic;
SIGNAL N2_74 : std_logic;
SIGNAL N2_75 : std_logic;
SIGNAL N2_76 : std_logic;
SIGNAL N2_77 : std_logic;
SIGNAL N2_78 : std_logic;
SIGNAL N2_79 : std_logic;
SIGNAL N2_80 : std_logic;
SIGNAL N2_81 : std_logic;
SIGNAL N2_82 : std_logic;
SIGNAL N2_83 : std_logic;
SIGNAL N2_84 : std_logic;
SIGNAL N2_85 : std_logic;
SIGNAL N3_0 : std_logic;
SIGNAL N3_1 : std_logic;
SIGNAL N3_2 : std_logic;
SIGNAL N3_3 : std_logic;
SIGNAL N3_4 : std_logic;
SIGNAL N3_5 : std_logic;
SIGNAL N3_6 : std_logic;
SIGNAL N3_7 : std_logic;
SIGNAL N3_8 : std_logic;
SIGNAL N3_9 : std_logic;
SIGNAL N3_10 : std_logic;
SIGNAL N3_11 : std_logic;
SIGNAL N3_12 : std_logic;
SIGNAL N3_13 : std_logic;
SIGNAL N3_14 : std_logic;
SIGNAL H3_0 : std_logic;
SIGNAL C3_0 : std_logic;
SIGNAL N3_15 : std_logic;
SIGNAL N3_16 : std_logic;
SIGNAL N3_17 : std_logic;
SIGNAL H3_1 : std_logic;
SIGNAL C3_1 : std_logic;
SIGNAL N3_18 : std_logic;
SIGNAL N3_19 : std_logic;
SIGNAL F3_0 : std_logic;
SIGNAL C3_2 : std_logic;
SIGNAL H3_2 : std_logic;
SIGNAL C3_3 : std_logic;
SIGNAL N3_20 : std_logic;
SIGNAL F3_1 : std_logic;
SIGNAL C3_4 : std_logic;
SIGNAL H3_3 : std_logic;
SIGNAL C3_5 : std_logic;
SIGNAL F3_2 : std_logic;
SIGNAL C3_6 : std_logic;
SIGNAL F3_3 : std_logic;
SIGNAL C3_7 : std_logic;
SIGNAL F3_4 : std_logic;
SIGNAL C3_8 : std_logic;
SIGNAL F3_5 : std_logic;
SIGNAL C3_9 : std_logic;
SIGNAL F3_6 : std_logic;
SIGNAL C3_10 : std_logic;
SIGNAL F3_7 : std_logic;
SIGNAL C3_11 : std_logic;
SIGNAL F3_8 : std_logic;
SIGNAL C3_12 : std_logic;
SIGNAL F3_9 : std_logic;
SIGNAL C3_13 : std_logic;
SIGNAL F3_10 : std_logic;
SIGNAL C3_14 : std_logic;
SIGNAL F3_11 : std_logic;
SIGNAL C3_15 : std_logic;
SIGNAL F3_12 : std_logic;
SIGNAL C3_16 : std_logic;
SIGNAL F3_13 : std_logic;
SIGNAL C3_17 : std_logic;
SIGNAL F3_14 : std_logic;
SIGNAL C3_18 : std_logic;
SIGNAL F3_15 : std_logic;
SIGNAL C3_19 : std_logic;
SIGNAL F3_16 : std_logic;
SIGNAL C3_20 : std_logic;
SIGNAL F3_17 : std_logic;
SIGNAL C3_21 : std_logic;
SIGNAL F3_18 : std_logic;
SIGNAL C3_22 : std_logic;
SIGNAL F3_19 : std_logic;
SIGNAL C3_23 : std_logic;
SIGNAL F3_20 : std_logic;
SIGNAL C3_24 : std_logic;
SIGNAL F3_21 : std_logic;
SIGNAL C3_25 : std_logic;
SIGNAL F3_22 : std_logic;
SIGNAL C3_26 : std_logic;
SIGNAL F3_23 : std_logic;
SIGNAL C3_27 : std_logic;
SIGNAL F3_24 : std_logic;
SIGNAL C3_28 : std_logic;
SIGNAL F3_25 : std_logic;
SIGNAL C3_29 : std_logic;
SIGNAL F3_26 : std_logic;
SIGNAL C3_30 : std_logic;
SIGNAL F3_27 : std_logic;
SIGNAL C3_31 : std_logic;
SIGNAL F3_28 : std_logic;
SIGNAL C3_32 : std_logic;
SIGNAL F3_29 : std_logic;
SIGNAL C3_33 : std_logic;
SIGNAL F3_30 : std_logic;
SIGNAL C3_34 : std_logic;
SIGNAL F3_31 : std_logic;
SIGNAL C3_35 : std_logic;
SIGNAL F3_32 : std_logic;
SIGNAL C3_36 : std_logic;
SIGNAL F3_33 : std_logic;
SIGNAL C3_37 : std_logic;
SIGNAL F3_34 : std_logic;
SIGNAL C3_38 : std_logic;
SIGNAL F3_35 : std_logic;
SIGNAL C3_39 : std_logic;
SIGNAL F3_36 : std_logic;
SIGNAL C3_40 : std_logic;
SIGNAL F3_37 : std_logic;
SIGNAL C3_41 : std_logic;
SIGNAL F3_38 : std_logic;
SIGNAL C3_42 : std_logic;
SIGNAL F3_39 : std_logic;
SIGNAL C3_43 : std_logic;
SIGNAL F3_40 : std_logic;
SIGNAL C3_44 : std_logic;
SIGNAL F3_41 : std_logic;
SIGNAL C3_45 : std_logic;
SIGNAL F3_42 : std_logic;
SIGNAL C3_46 : std_logic;
SIGNAL F3_43 : std_logic;
SIGNAL C3_47 : std_logic;
SIGNAL F3_44 : std_logic;
SIGNAL C3_48 : std_logic;
SIGNAL F3_45 : std_logic;
SIGNAL C3_49 : std_logic;
SIGNAL F3_46 : std_logic;
SIGNAL C3_50 : std_logic;
SIGNAL F3_47 : std_logic;
SIGNAL C3_51 : std_logic;
SIGNAL F3_48 : std_logic;
SIGNAL C3_52 : std_logic;
SIGNAL F3_49 : std_logic;
SIGNAL C3_53 : std_logic;
SIGNAL F3_50 : std_logic;
SIGNAL C3_54 : std_logic;
SIGNAL F3_51 : std_logic;
SIGNAL C3_55 : std_logic;
SIGNAL F3_52 : std_logic;
SIGNAL C3_56 : std_logic;
SIGNAL F3_53 : std_logic;
SIGNAL C3_57 : std_logic;
SIGNAL F3_54 : std_logic;
SIGNAL C3_58 : std_logic;
SIGNAL F3_55 : std_logic;
SIGNAL C3_59 : std_logic;
SIGNAL F3_56 : std_logic;
SIGNAL C3_60 : std_logic;
SIGNAL F3_57 : std_logic;
SIGNAL C3_61 : std_logic;
SIGNAL F3_58 : std_logic;
SIGNAL C3_62 : std_logic;
SIGNAL F3_59 : std_logic;
SIGNAL C3_63 : std_logic;
SIGNAL F3_60 : std_logic;
SIGNAL C3_64 : std_logic;
SIGNAL F3_61 : std_logic;
SIGNAL C3_65 : std_logic;
SIGNAL F3_62 : std_logic;
SIGNAL C3_66 : std_logic;
SIGNAL F3_63 : std_logic;
SIGNAL C3_67 : std_logic;
SIGNAL F3_64 : std_logic;
SIGNAL C3_68 : std_logic;
SIGNAL F3_65 : std_logic;
SIGNAL C3_69 : std_logic;
SIGNAL F3_66 : std_logic;
SIGNAL C3_70 : std_logic;
SIGNAL H3_4 : std_logic;
SIGNAL C3_71 : std_logic;
SIGNAL F3_67 : std_logic;
SIGNAL C3_72 : std_logic;
SIGNAL N3_21 : std_logic;
SIGNAL H3_5 : std_logic;
SIGNAL C3_73 : std_logic;
SIGNAL N3_22 : std_logic;
SIGNAL N3_23 : std_logic;
SIGNAL N3_24 : std_logic;
SIGNAL N3_25 : std_logic;
SIGNAL N3_26 : std_logic;
SIGNAL N3_27 : std_logic;
SIGNAL N3_28 : std_logic;
SIGNAL N3_29 : std_logic;
SIGNAL N3_30 : std_logic;
SIGNAL N3_31 : std_logic;
SIGNAL N4_0 : std_logic;
SIGNAL N4_1 : std_logic;
SIGNAL N4_2 : std_logic;
SIGNAL N4_3 : std_logic;
SIGNAL N4_4 : std_logic;
SIGNAL N4_5 : std_logic;
SIGNAL N4_6 : std_logic;
SIGNAL N4_7 : std_logic;
SIGNAL H4_0 : std_logic;
SIGNAL C4_0 : std_logic;
SIGNAL N4_8 : std_logic;
SIGNAL N4_9 : std_logic;
SIGNAL H4_1 : std_logic;
SIGNAL C4_1 : std_logic;
SIGNAL N4_10 : std_logic;
SIGNAL F4_0 : std_logic;
SIGNAL C4_2 : std_logic;
SIGNAL N4_11 : std_logic;
SIGNAL F4_1 : std_logic;
SIGNAL C4_3 : std_logic;
SIGNAL N4_12 : std_logic;
SIGNAL F4_2 : std_logic;
SIGNAL C4_4 : std_logic;
SIGNAL N4_13 : std_logic;
SIGNAL F4_3 : std_logic;
SIGNAL C4_5 : std_logic;
SIGNAL N4_14 : std_logic;
SIGNAL F4_4 : std_logic;
SIGNAL C4_6 : std_logic;
SIGNAL N4_15 : std_logic;
SIGNAL F4_5 : std_logic;
SIGNAL C4_7 : std_logic;
SIGNAL N4_16 : std_logic;
SIGNAL F4_6 : std_logic;
SIGNAL C4_8 : std_logic;
SIGNAL N4_17 : std_logic;
SIGNAL F4_7 : std_logic;
SIGNAL C4_9 : std_logic;
SIGNAL N4_18 : std_logic;
SIGNAL F4_8 : std_logic;
SIGNAL C4_10 : std_logic;
SIGNAL N4_19 : std_logic;
SIGNAL F4_9 : std_logic;
SIGNAL C4_11 : std_logic;
SIGNAL N4_20 : std_logic;
SIGNAL F4_10 : std_logic;
SIGNAL C4_12 : std_logic;
SIGNAL N4_21 : std_logic;
SIGNAL F4_11 : std_logic;
SIGNAL C4_13 : std_logic;
SIGNAL N4_22 : std_logic;
SIGNAL F4_12 : std_logic;
SIGNAL C4_14 : std_logic;
SIGNAL N4_23 : std_logic;
SIGNAL F4_13 : std_logic;
SIGNAL C4_15 : std_logic;
SIGNAL N4_24 : std_logic;
SIGNAL F4_14 : std_logic;
SIGNAL C4_16 : std_logic;
SIGNAL N4_25 : std_logic;
SIGNAL F4_15 : std_logic;
SIGNAL C4_17 : std_logic;
SIGNAL N4_26 : std_logic;
SIGNAL F4_16 : std_logic;
SIGNAL C4_18 : std_logic;
SIGNAL N4_27 : std_logic;
SIGNAL F4_17 : std_logic;
SIGNAL C4_19 : std_logic;
SIGNAL N4_28 : std_logic;
SIGNAL F4_18 : std_logic;
SIGNAL C4_20 : std_logic;
SIGNAL N4_29 : std_logic;
SIGNAL F4_19 : std_logic;
SIGNAL C4_21 : std_logic;
SIGNAL N4_30 : std_logic;
SIGNAL F4_20 : std_logic;
SIGNAL C4_22 : std_logic;
SIGNAL N4_31 : std_logic;
SIGNAL F4_21 : std_logic;
SIGNAL C4_23 : std_logic;
SIGNAL N4_32 : std_logic;
SIGNAL F4_22 : std_logic;
SIGNAL C4_24 : std_logic;
SIGNAL N4_33 : std_logic;
SIGNAL F4_23 : std_logic;
SIGNAL C4_25 : std_logic;
SIGNAL N4_34 : std_logic;
SIGNAL F4_24 : std_logic;
SIGNAL C4_26 : std_logic;
SIGNAL N4_35 : std_logic;
SIGNAL F4_25 : std_logic;
SIGNAL C4_27 : std_logic;
SIGNAL N4_36 : std_logic;
SIGNAL F4_26 : std_logic;
SIGNAL C4_28 : std_logic;
SIGNAL N4_37 : std_logic;
SIGNAL F4_27 : std_logic;
SIGNAL C4_29 : std_logic;
SIGNAL N4_38 : std_logic;
SIGNAL F4_28 : std_logic;
SIGNAL C4_30 : std_logic;
SIGNAL N4_39 : std_logic;
SIGNAL F4_29 : std_logic;
SIGNAL C4_31 : std_logic;
SIGNAL N4_40 : std_logic;
SIGNAL F4_30 : std_logic;
SIGNAL C4_32 : std_logic;
SIGNAL N4_41 : std_logic;
SIGNAL F4_31 : std_logic;
SIGNAL C4_33 : std_logic;
SIGNAL N4_42 : std_logic;
SIGNAL F4_32 : std_logic;
SIGNAL C4_34 : std_logic;
SIGNAL N4_43 : std_logic;
SIGNAL F4_33 : std_logic;
SIGNAL C4_35 : std_logic;
SIGNAL N4_44 : std_logic;
SIGNAL F4_34 : std_logic;
SIGNAL C4_36 : std_logic;
SIGNAL N4_45 : std_logic;
SIGNAL F4_35 : std_logic;
SIGNAL C4_37 : std_logic;
SIGNAL N4_46 : std_logic;
SIGNAL F4_36 : std_logic;
SIGNAL C4_38 : std_logic;
SIGNAL N4_47 : std_logic;
SIGNAL F4_37 : std_logic;
SIGNAL C4_39 : std_logic;
SIGNAL N4_48 : std_logic;
SIGNAL F4_38 : std_logic;
SIGNAL C4_40 : std_logic;
SIGNAL N4_49 : std_logic;
SIGNAL F4_39 : std_logic;
SIGNAL C4_41 : std_logic;
SIGNAL N4_50 : std_logic;
SIGNAL H4_2 : std_logic;
SIGNAL C4_42 : std_logic;
SIGNAL N4_51 : std_logic;
SIGNAL N4_52 : std_logic;
SIGNAL N4_53 : std_logic;
SIGNAL N5_0 : std_logic;
SIGNAL N5_1 : std_logic;
SIGNAL N5_2 : std_logic;
SIGNAL H5_0 : std_logic;
SIGNAL C5_0 : std_logic;
SIGNAL N5_3 : std_logic;
SIGNAL H5_1 : std_logic;
SIGNAL C5_1 : std_logic;
SIGNAL F5_0 : std_logic;
SIGNAL C5_2 : std_logic;
SIGNAL F5_1 : std_logic;
SIGNAL C5_3 : std_logic;
SIGNAL F5_2 : std_logic;
SIGNAL C5_4 : std_logic;
SIGNAL F5_3 : std_logic;
SIGNAL C5_5 : std_logic;
SIGNAL F5_4 : std_logic;
SIGNAL C5_6 : std_logic;
SIGNAL F5_5 : std_logic;
SIGNAL C5_7 : std_logic;
SIGNAL F5_6 : std_logic;
SIGNAL C5_8 : std_logic;
SIGNAL F5_7 : std_logic;
SIGNAL C5_9 : std_logic;
SIGNAL F5_8 : std_logic;
SIGNAL C5_10 : std_logic;
SIGNAL F5_9 : std_logic;
SIGNAL C5_11 : std_logic;
SIGNAL F5_10 : std_logic;
SIGNAL C5_12 : std_logic;
SIGNAL F5_11 : std_logic;
SIGNAL C5_13 : std_logic;
SIGNAL F5_12 : std_logic;
SIGNAL C5_14 : std_logic;
SIGNAL F5_13 : std_logic;
SIGNAL C5_15 : std_logic;
SIGNAL F5_14 : std_logic;
SIGNAL C5_16 : std_logic;
SIGNAL F5_15 : std_logic;
SIGNAL C5_17 : std_logic;
SIGNAL F5_16 : std_logic;
SIGNAL C5_18 : std_logic;
SIGNAL F5_17 : std_logic;
SIGNAL C5_19 : std_logic;
SIGNAL F5_18 : std_logic;
SIGNAL C5_20 : std_logic;
SIGNAL F5_19 : std_logic;
SIGNAL C5_21 : std_logic;
SIGNAL F5_20 : std_logic;
SIGNAL C5_22 : std_logic;
SIGNAL F5_21 : std_logic;
SIGNAL C5_23 : std_logic;
SIGNAL F5_22 : std_logic;
SIGNAL C5_24 : std_logic;
SIGNAL F5_23 : std_logic;
SIGNAL C5_25 : std_logic;
SIGNAL F5_24 : std_logic;
SIGNAL C5_26 : std_logic;
SIGNAL F5_25 : std_logic;
SIGNAL C5_27 : std_logic;
SIGNAL F5_26 : std_logic;
SIGNAL C5_28 : std_logic;
SIGNAL F5_27 : std_logic;
SIGNAL C5_29 : std_logic;
SIGNAL F5_28 : std_logic;
SIGNAL C5_30 : std_logic;
SIGNAL F5_29 : std_logic;
SIGNAL C5_31 : std_logic;
SIGNAL F5_30 : std_logic;
SIGNAL C5_32 : std_logic;
SIGNAL F5_31 : std_logic;
SIGNAL C5_33 : std_logic;
SIGNAL F5_32 : std_logic;
SIGNAL C5_34 : std_logic;
SIGNAL F5_33 : std_logic;
SIGNAL C5_35 : std_logic;
SIGNAL F5_34 : std_logic;
SIGNAL C5_36 : std_logic;
SIGNAL F5_35 : std_logic;
SIGNAL C5_37 : std_logic;
SIGNAL F5_36 : std_logic;
SIGNAL C5_38 : std_logic;
SIGNAL F5_37 : std_logic;
SIGNAL C5_39 : std_logic;
SIGNAL F5_38 : std_logic;
SIGNAL C5_40 : std_logic;
SIGNAL F5_39 : std_logic;
SIGNAL C5_41 : std_logic;
SIGNAL F5_40 : std_logic;
SIGNAL C5_42 : std_logic;
SIGNAL F5_41 : std_logic;
SIGNAL C5_43 : std_logic;
SIGNAL F5_42 : std_logic;
SIGNAL C5_44 : std_logic;
SIGNAL F5_43 : std_logic;
SIGNAL Co_0 : std_logic;
SIGNAL Co_1 : std_logic;
SIGNAL Co_2 : std_logic;
SIGNAL Co_3 : std_logic;
SIGNAL Co_4 : std_logic;
SIGNAL Co_5 : std_logic;
SIGNAL Co_6 : std_logic;
SIGNAL Co_7 : std_logic;
SIGNAL Co_8 : std_logic;
SIGNAL Co_9 : std_logic;
SIGNAL Co_10 : std_logic;
SIGNAL Co_11 : std_logic;
SIGNAL Co_12 : std_logic;
SIGNAL Co_13 : std_logic;
SIGNAL Co_14 : std_logic;
SIGNAL Co_15 : std_logic;
SIGNAL Co_16 : std_logic;
SIGNAL Co_17 : std_logic;
SIGNAL Co_18 : std_logic;
SIGNAL Co_19 : std_logic;
SIGNAL Co_20 : std_logic;
SIGNAL Co_21 : std_logic;
SIGNAL Co_22 : std_logic;
SIGNAL Co_23 : std_logic;
SIGNAL Co_24 : std_logic;
SIGNAL Co_25 : std_logic;
SIGNAL Co_26 : std_logic;
SIGNAL Co_27 : std_logic;
SIGNAL Co_28 : std_logic;
SIGNAL Co_29 : std_logic;
SIGNAL Co_30 : std_logic;
SIGNAL Co_31 : std_logic;
SIGNAL Co_32 : std_logic;
SIGNAL Co_33 : std_logic;
SIGNAL Co_34 : std_logic;
SIGNAL Co_35 : std_logic;
SIGNAL Co_36 : std_logic;
SIGNAL Co_37 : std_logic;
SIGNAL Co_38 : std_logic;
SIGNAL Co_39 : std_logic;
SIGNAL Co_40 : std_logic;
SIGNAL Co_41 : std_logic;
SIGNAL Co_42 : std_logic;
SIGNAL Co_43 : std_logic;
SIGNAL Co_44 : std_logic;
SIGNAL Co_45 : std_logic;
SIGNAL Co_46 : std_logic;

COMPONENT FA IS
PORT(I1 : IN std_logic;
I2 : IN std_logic;
Cin : IN std_logic;
Q : OUT std_logic;
Cout : OUT std_logic);
END COMPONENT;

COMPONENT HA IS
PORT(I1 : IN std_logic;
I2 : IN std_logic;
Q : OUT std_logic;
Cout : OUT std_logic);
END COMPONENT;

BEGIN

N0_358 <= Li(26);
N0_359 <= Mi(24);
N0_355 <= Ki(27);
N0_356 <= Li(25);
N0_357 <= Mi(23);
N0_352 <= Ki(26);
N0_353 <= Li(24);
N0_354 <= Mi(22);
N0_348 <= Ji(27);
N0_349 <= Ki(25);
N0_350 <= Li(23);
N0_351 <= Mi(21);
N0_344 <= Ji(26);
N0_345 <= Ki(24);
N0_346 <= Li(22);
N0_347 <= Mi(20);
N0_339 <= Ii(27);
N0_340 <= Ji(25);
N0_341 <= Ki(23);
N0_342 <= Li(21);
N0_343 <= Mi(19);
N0_334 <= Ii(26);
N0_335 <= Ji(24);
N0_336 <= Ki(22);
N0_337 <= Li(20);
N0_338 <= Mi(18);
N0_328 <= Hi(27);
N0_329 <= Ii(25);
N0_330 <= Ji(23);
N0_331 <= Ki(21);
N0_332 <= Li(19);
N0_333 <= Mi(17);
N0_322 <= Hi(26);
N0_323 <= Ii(24);
N0_324 <= Ji(22);
N0_325 <= Ki(20);
N0_326 <= Li(18);
N0_327 <= Mi(16);
N0_315 <= Gi(27);
N0_316 <= Hi(25);
N0_317 <= Ii(23);
N0_318 <= Ji(21);
N0_319 <= Ki(19);
N0_320 <= Li(17);
N0_321 <= Mi(15);
N0_308 <= Gi(26);
N0_309 <= Hi(24);
N0_310 <= Ii(22);
N0_311 <= Ji(20);
N0_312 <= Ki(18);
N0_313 <= Li(16);
N0_314 <= Mi(14);
N0_300 <= Fi(27);
N0_301 <= Gi(25);
N0_302 <= Hi(23);
N0_303 <= Ii(21);
N0_304 <= Ji(19);
N0_305 <= Ki(17);
N0_306 <= Li(15);
N0_307 <= Mi(13);
N0_292 <= Fi(26);
N0_293 <= Gi(24);
N0_294 <= Hi(22);
N0_295 <= Ii(20);
N0_296 <= Ji(18);
N0_297 <= Ki(16);
N0_298 <= Li(14);
N0_299 <= Mi(12);
N0_283 <= Ei(27);
N0_284 <= Fi(25);
N0_285 <= Gi(23);
N0_286 <= Hi(21);
N0_287 <= Ii(19);
N0_288 <= Ji(17);
N0_289 <= Ki(15);
N0_290 <= Li(13);
N0_291 <= Mi(11);
N0_274 <= Ei(26);
N0_275 <= Fi(24);
N0_276 <= Gi(22);
N0_277 <= Hi(20);
N0_278 <= Ii(18);
N0_279 <= Ji(16);
N0_280 <= Ki(14);
N0_281 <= Li(12);
N0_282 <= Mi(10);
N0_264 <= Di(27);
N0_265 <= Ei(25);
N0_266 <= Fi(23);
N0_267 <= Gi(21);
N0_268 <= Hi(19);
N0_269 <= Ii(17);
N0_270 <= Ji(15);
N0_271 <= Ki(13);
N0_272 <= Li(11);
N0_273 <= Mi(9);
N0_254 <= Di(26);
N0_255 <= Ei(24);
N0_256 <= Fi(22);
N0_257 <= Gi(20);
N0_258 <= Hi(18);
N0_259 <= Ii(16);
N0_260 <= Ji(14);
N0_261 <= Ki(12);
N0_262 <= Li(10);
N0_263 <= Mi(8);
N0_243 <= Ci(27);
N0_244 <= Di(25);
N0_245 <= Ei(23);
N0_246 <= Fi(21);
N0_247 <= Gi(19);
N0_248 <= Hi(17);
N0_249 <= Ii(15);
N0_250 <= Ji(13);
N0_251 <= Ki(11);
N0_252 <= Li(9);
N0_253 <= Mi(7);
N0_232 <= Ci(26);
N0_233 <= Di(24);
N0_234 <= Ei(22);
N0_235 <= Fi(20);
N0_236 <= Gi(18);
N0_237 <= Hi(16);
N0_238 <= Ii(14);
N0_239 <= Ji(12);
N0_240 <= Ki(10);
N0_241 <= Li(8);
N0_242 <= Mi(6);
N0_220 <= Bi(27);
N0_221 <= Ci(25);
N0_222 <= Di(23);
N0_223 <= Ei(21);
N0_224 <= Fi(19);
N0_225 <= Gi(17);
N0_226 <= Hi(15);
N0_227 <= Ii(13);
N0_228 <= Ji(11);
N0_229 <= Ki(9);
N0_230 <= Li(7);
N0_231 <= Mi(5);
N0_207 <= Ai(27);
N0_208 <= Bi(26);
N0_209 <= Ci(24);
N0_210 <= Di(22);
N0_211 <= Ei(20);
N0_212 <= Fi(18);
N0_213 <= Gi(16);
N0_214 <= Hi(14);
N0_215 <= Ii(12);
N0_216 <= Ji(10);
N0_217 <= Ki(8);
N0_218 <= Li(6);
N0_219 <= Mi(4);
N0_194 <= Ai(26);
N0_195 <= Bi(25);
N0_196 <= Ci(23);
N0_197 <= Di(21);
N0_198 <= Ei(19);
N0_199 <= Fi(17);
N0_200 <= Gi(15);
N0_201 <= Hi(13);
N0_202 <= Ii(11);
N0_203 <= Ji(9);
N0_204 <= Ki(7);
N0_205 <= Li(5);
N0_206 <= Mi(3);
N0_181 <= Ai(25);
N0_182 <= Bi(24);
N0_183 <= Ci(22);
N0_184 <= Di(20);
N0_185 <= Ei(18);
N0_186 <= Fi(16);
N0_187 <= Gi(14);
N0_188 <= Hi(12);
N0_189 <= Ii(10);
N0_190 <= Ji(8);
N0_191 <= Ki(6);
N0_192 <= Li(4);
N0_193 <= Mi(2);
N0_168 <= Ai(24);
N0_169 <= Bi(23);
N0_170 <= Ci(21);
N0_171 <= Di(19);
N0_172 <= Ei(17);
N0_173 <= Fi(15);
N0_174 <= Gi(13);
N0_175 <= Hi(11);
N0_176 <= Ii(9);
N0_177 <= Ji(7);
N0_178 <= Ki(5);
N0_179 <= Li(3);
N0_180 <= Mi(1);
N0_156 <= Ai(23);
N0_157 <= Bi(22);
N0_158 <= Ci(20);
N0_159 <= Di(18);
N0_160 <= Ei(16);
N0_161 <= Fi(14);
N0_162 <= Gi(12);
N0_163 <= Hi(10);
N0_164 <= Ii(8);
N0_165 <= Ji(6);
N0_166 <= Ki(4);
N0_167 <= Li(2);
N0_143 <= Ai(22);
N0_144 <= Bi(21);
N0_145 <= Ci(19);
N0_146 <= Di(17);
N0_147 <= Ei(15);
N0_148 <= Fi(13);
N0_149 <= Gi(11);
N0_150 <= Hi(9);
N0_151 <= Ii(7);
N0_152 <= Ji(5);
N0_153 <= Ki(3);
N0_154 <= Li(1);
N0_155 <= Mi(0);
N0_132 <= Ai(21);
N0_133 <= Bi(20);
N0_134 <= Ci(18);
N0_135 <= Di(16);
N0_136 <= Ei(14);
N0_137 <= Fi(12);
N0_138 <= Gi(10);
N0_139 <= Hi(8);
N0_140 <= Ii(6);
N0_141 <= Ji(4);
N0_142 <= Ki(2);
N0_120 <= Ai(20);
N0_121 <= Bi(19);
N0_122 <= Ci(17);
N0_123 <= Di(15);
N0_124 <= Ei(13);
N0_125 <= Fi(11);
N0_126 <= Gi(9);
N0_127 <= Hi(7);
N0_128 <= Ii(5);
N0_129 <= Ji(3);
N0_130 <= Ki(1);
N0_131 <= Li(0);
N0_110 <= Ai(19);
N0_111 <= Bi(18);
N0_112 <= Ci(16);
N0_113 <= Di(14);
N0_114 <= Ei(12);
N0_115 <= Fi(10);
N0_116 <= Gi(8);
N0_117 <= Hi(6);
N0_118 <= Ii(4);
N0_119 <= Ji(2);
N0_99 <= Ai(18);
N0_100 <= Bi(17);
N0_101 <= Ci(15);
N0_102 <= Di(13);
N0_103 <= Ei(11);
N0_104 <= Fi(9);
N0_105 <= Gi(7);
N0_106 <= Hi(5);
N0_107 <= Ii(3);
N0_108 <= Ji(1);
N0_109 <= Ki(0);
N0_90 <= Ai(17);
N0_91 <= Bi(16);
N0_92 <= Ci(14);
N0_93 <= Di(12);
N0_94 <= Ei(10);
N0_95 <= Fi(8);
N0_96 <= Gi(6);
N0_97 <= Hi(4);
N0_98 <= Ii(2);
N0_80 <= Ai(16);
N0_81 <= Bi(15);
N0_82 <= Ci(13);
N0_83 <= Di(11);
N0_84 <= Ei(9);
N0_85 <= Fi(7);
N0_86 <= Gi(5);
N0_87 <= Hi(3);
N0_88 <= Ii(1);
N0_89 <= Ji(0);
N0_72 <= Ai(15);
N0_73 <= Bi(14);
N0_74 <= Ci(12);
N0_75 <= Di(10);
N0_76 <= Ei(8);
N0_77 <= Fi(6);
N0_78 <= Gi(4);
N0_79 <= Hi(2);
N0_63 <= Ai(14);
N0_64 <= Bi(13);
N0_65 <= Ci(11);
N0_66 <= Di(9);
N0_67 <= Ei(7);
N0_68 <= Fi(5);
N0_69 <= Gi(3);
N0_70 <= Hi(1);
N0_71 <= Ii(0);
N0_56 <= Ai(13);
N0_57 <= Bi(12);
N0_58 <= Ci(10);
N0_59 <= Di(8);
N0_60 <= Ei(6);
N0_61 <= Fi(4);
N0_62 <= Gi(2);
N0_48 <= Ai(12);
N0_49 <= Bi(11);
N0_50 <= Ci(9);
N0_51 <= Di(7);
N0_52 <= Ei(5);
N0_53 <= Fi(3);
N0_54 <= Gi(1);
N0_55 <= Hi(0);
N0_42 <= Ai(11);
N0_43 <= Bi(10);
N0_44 <= Ci(8);
N0_45 <= Di(6);
N0_46 <= Ei(4);
N0_47 <= Fi(2);
N0_35 <= Ai(10);
N0_36 <= Bi(9);
N0_37 <= Ci(7);
N0_38 <= Di(5);
N0_39 <= Ei(3);
N0_40 <= Fi(1);
N0_41 <= Gi(0);
N0_30 <= Ai(9);
N0_31 <= Bi(8);
N0_32 <= Ci(6);
N0_33 <= Di(4);
N0_34 <= Ei(2);
N0_24 <= Ai(8);
N0_25 <= Bi(7);
N0_26 <= Ci(5);
N0_27 <= Di(3);
N0_28 <= Ei(1);
N0_29 <= Fi(0);
N0_20 <= Ai(7);
N0_21 <= Bi(6);
N0_22 <= Ci(4);
N0_23 <= Di(2);
N0_15 <= Ai(6);
N0_16 <= Bi(5);
N0_17 <= Ci(3);
N0_18 <= Di(1);
N0_19 <= Ei(0);
N0_12 <= Ai(5);
N0_13 <= Bi(4);
N0_14 <= Ci(2);
N0_8 <= Ai(4);
N0_9 <= Bi(3);
N0_10 <= Ci(1);
N0_11 <= Di(0);
N0_6 <= Ai(3);
N0_7 <= Bi(2);
N0_3 <= Ai(2);
N0_4 <= Bi(1);
N0_5 <= Ci(0);
N0_2 <= Ai(1);
N0_0 <= Ai(0);
N0_1 <= Bi(0);
N1_0 <= N0_0;
N1_1 <= N0_1;
N1_2 <= N0_2;
N1_3 <= N0_3;
N1_4 <= N0_4;
N1_5 <= N0_5;
N1_6 <= N0_6;
N1_7 <= N0_7;
N1_8 <= N0_8;
N1_9 <= N0_9;
N1_10 <= N0_10;
N1_11 <= N0_11;
N1_12 <= N0_12;
N1_13 <= N0_13;
N1_14 <= N0_14;
N1_15 <= N0_15;
N1_16 <= N0_16;
N1_17 <= N0_17;
N1_18 <= N0_18;
N1_19 <= N0_19;
N1_20 <= N0_20;
N1_21 <= N0_21;
N1_22 <= N0_22;
N1_23 <= N0_23;
N1_24 <= N0_24;
N1_25 <= N0_25;
N1_26 <= N0_26;
N1_27 <= N0_27;
N1_28 <= N0_28;
N1_29 <= N0_29;
N1_30 <= N0_30;
N1_31 <= N0_31;
N1_32 <= N0_32;
N1_33 <= N0_33;
N1_34 <= N0_34;
N1_35 <= N0_35;
N1_36 <= N0_36;
N1_37 <= N0_37;
N1_38 <= N0_38;
N1_39 <= N0_39;
N1_40 <= N0_40;
N1_41 <= N0_41;
N1_42 <= N0_42;
N1_43 <= N0_43;
N1_44 <= N0_44;
N1_45 <= N0_45;
N1_46 <= N0_46;
N1_47 <= N0_47;
N1_48 <= N0_48;
N1_49 <= N0_49;
N1_50 <= N0_50;
N1_51 <= N0_51;
N1_52 <= N0_52;
N1_53 <= N0_53;
N1_54 <= N0_54;
N1_55 <= N0_55;
N1_56 <= N0_56;
N1_57 <= N0_57;
N1_58 <= N0_58;
N1_59 <= N0_59;
N1_60 <= N0_60;
N1_61 <= N0_61;
N1_62 <= N0_62;
N1_63 <= N0_63;
N1_64 <= N0_64;
N1_65 <= N0_65;
N1_66 <= N0_66;
N1_67 <= N0_67;
N1_68 <= N0_68;
N1_69 <= N0_69;
N1_70 <= N0_70;
N1_71 <= N0_71;
N1_72 <= N0_72;
N1_73 <= N0_73;
N1_74 <= N0_74;
N1_75 <= N0_75;
N1_76 <= N0_76;
N1_77 <= N0_77;
N1_78 <= N0_78;
N1_79 <= N0_79;
H0 : HA PORT MAP(N0_80,N0_81,H1_0,C1_0);
N1_80 <= N0_82;
N1_81 <= N0_83;
N1_82 <= N0_84;
N1_83 <= N0_85;
N1_84 <= N0_86;
N1_85 <= N0_87;
N1_86 <= N0_88;
N1_87 <= N0_89;
H1 : HA PORT MAP(N0_90,N0_91,H1_1,C1_1);
N1_88 <= N0_92;
N1_89 <= N0_93;
N1_90 <= N0_94;
N1_91 <= N0_95;
N1_92 <= N0_96;
N1_93 <= N0_97;
N1_94 <= N0_98;
F0 : FA PORT MAP(N0_99,N0_100,N0_101,F1_0,C1_2);
H2 : HA PORT MAP(N0_102,N0_103,H1_2,C1_3);
N1_95 <= N0_104;
N1_96 <= N0_105;
N1_97 <= N0_106;
N1_98 <= N0_107;
N1_99 <= N0_108;
N1_100 <= N0_109;
F1 : FA PORT MAP(N0_110,N0_111,N0_112,F1_1,C1_4);
H3 : HA PORT MAP(N0_113,N0_114,H1_3,C1_5);
N1_101 <= N0_115;
N1_102 <= N0_116;
N1_103 <= N0_117;
N1_104 <= N0_118;
N1_105 <= N0_119;
F2 : FA PORT MAP(N0_120,N0_121,N0_122,F1_2,C1_6);
F3 : FA PORT MAP(N0_123,N0_124,N0_125,F1_3,C1_7);
H4 : HA PORT MAP(N0_126,N0_127,H1_4,C1_8);
N1_106 <= N0_128;
N1_107 <= N0_129;
N1_108 <= N0_130;
N1_109 <= N0_131;
F4 : FA PORT MAP(N0_132,N0_133,N0_134,F1_4,C1_9);
F5 : FA PORT MAP(N0_135,N0_136,N0_137,F1_5,C1_10);
H5 : HA PORT MAP(N0_138,N0_139,H1_5,C1_11);
N1_110 <= N0_140;
N1_111 <= N0_141;
N1_112 <= N0_142;
F6 : FA PORT MAP(N0_143,N0_144,N0_145,F1_6,C1_12);
F7 : FA PORT MAP(N0_146,N0_147,N0_148,F1_7,C1_13);
F8 : FA PORT MAP(N0_149,N0_150,N0_151,F1_8,C1_14);
H6 : HA PORT MAP(N0_152,N0_153,H1_6,C1_15);
N1_113 <= N0_154;
N1_114 <= N0_155;
F9 : FA PORT MAP(N0_156,N0_157,N0_158,F1_9,C1_16);
F10 : FA PORT MAP(N0_159,N0_160,N0_161,F1_10,C1_17);
F11 : FA PORT MAP(N0_162,N0_163,N0_164,F1_11,C1_18);
H7 : HA PORT MAP(N0_165,N0_166,H1_7,C1_19);
N1_115 <= N0_167;
F12 : FA PORT MAP(N0_168,N0_169,N0_170,F1_12,C1_20);
F13 : FA PORT MAP(N0_171,N0_172,N0_173,F1_13,C1_21);
F14 : FA PORT MAP(N0_174,N0_175,N0_176,F1_14,C1_22);
F15 : FA PORT MAP(N0_177,N0_178,N0_179,F1_15,C1_23);
N1_116 <= N0_180;
F16 : FA PORT MAP(N0_181,N0_182,N0_183,F1_16,C1_24);
F17 : FA PORT MAP(N0_184,N0_185,N0_186,F1_17,C1_25);
F18 : FA PORT MAP(N0_187,N0_188,N0_189,F1_18,C1_26);
F19 : FA PORT MAP(N0_190,N0_191,N0_192,F1_19,C1_27);
N1_117 <= N0_193;
F20 : FA PORT MAP(N0_194,N0_195,N0_196,F1_20,C1_28);
F21 : FA PORT MAP(N0_197,N0_198,N0_199,F1_21,C1_29);
F22 : FA PORT MAP(N0_200,N0_201,N0_202,F1_22,C1_30);
F23 : FA PORT MAP(N0_203,N0_204,N0_205,F1_23,C1_31);
N1_118 <= N0_206;
F24 : FA PORT MAP(N0_207,N0_208,N0_209,F1_24,C1_32);
F25 : FA PORT MAP(N0_210,N0_211,N0_212,F1_25,C1_33);
F26 : FA PORT MAP(N0_213,N0_214,N0_215,F1_26,C1_34);
F27 : FA PORT MAP(N0_216,N0_217,N0_218,F1_27,C1_35);
N1_119 <= N0_219;
F28 : FA PORT MAP(N0_220,N0_221,N0_222,F1_28,C1_36);
F29 : FA PORT MAP(N0_223,N0_224,N0_225,F1_29,C1_37);
F30 : FA PORT MAP(N0_226,N0_227,N0_228,F1_30,C1_38);
H8 : HA PORT MAP(N0_229,N0_230,H1_8,C1_39);
N1_120 <= N0_231;
F31 : FA PORT MAP(N0_232,N0_233,N0_234,F1_31,C1_40);
F32 : FA PORT MAP(N0_235,N0_236,N0_237,F1_32,C1_41);
F33 : FA PORT MAP(N0_238,N0_239,N0_240,F1_33,C1_42);
N1_121 <= N0_241;
N1_122 <= N0_242;
F34 : FA PORT MAP(N0_243,N0_244,N0_245,F1_34,C1_43);
F35 : FA PORT MAP(N0_246,N0_247,N0_248,F1_35,C1_44);
H9 : HA PORT MAP(N0_249,N0_250,H1_9,C1_45);
N1_123 <= N0_251;
N1_124 <= N0_252;
N1_125 <= N0_253;
F36 : FA PORT MAP(N0_254,N0_255,N0_256,F1_36,C1_46);
F37 : FA PORT MAP(N0_257,N0_258,N0_259,F1_37,C1_47);
N1_126 <= N0_260;
N1_127 <= N0_261;
N1_128 <= N0_262;
N1_129 <= N0_263;
F38 : FA PORT MAP(N0_264,N0_265,N0_266,F1_38,C1_48);
H10 : HA PORT MAP(N0_267,N0_268,H1_10,C1_49);
N1_130 <= N0_269;
N1_131 <= N0_270;
N1_132 <= N0_271;
N1_133 <= N0_272;
N1_134 <= N0_273;
F39 : FA PORT MAP(N0_274,N0_275,N0_276,F1_39,C1_50);
N1_135 <= N0_277;
N1_136 <= N0_278;
N1_137 <= N0_279;
N1_138 <= N0_280;
N1_139 <= N0_281;
N1_140 <= N0_282;
H11 : HA PORT MAP(N0_283,N0_284,H1_11,C1_51);
N1_141 <= N0_285;
N1_142 <= N0_286;
N1_143 <= N0_287;
N1_144 <= N0_288;
N1_145 <= N0_289;
N1_146 <= N0_290;
N1_147 <= N0_291;
N1_148 <= N0_292;
N1_149 <= N0_293;
N1_150 <= N0_294;
N1_151 <= N0_295;
N1_152 <= N0_296;
N1_153 <= N0_297;
N1_154 <= N0_298;
N1_155 <= N0_299;
N1_156 <= N0_300;
N1_157 <= N0_301;
N1_158 <= N0_302;
N1_159 <= N0_303;
N1_160 <= N0_304;
N1_161 <= N0_305;
N1_162 <= N0_306;
N1_163 <= N0_307;
N1_164 <= N0_308;
N1_165 <= N0_309;
N1_166 <= N0_310;
N1_167 <= N0_311;
N1_168 <= N0_312;
N1_169 <= N0_313;
N1_170 <= N0_314;
N1_171 <= N0_315;
N1_172 <= N0_316;
N1_173 <= N0_317;
N1_174 <= N0_318;
N1_175 <= N0_319;
N1_176 <= N0_320;
N1_177 <= N0_321;
N1_178 <= N0_322;
N1_179 <= N0_323;
N1_180 <= N0_324;
N1_181 <= N0_325;
N1_182 <= N0_326;
N1_183 <= N0_327;
N1_184 <= N0_328;
N1_185 <= N0_329;
N1_186 <= N0_330;
N1_187 <= N0_331;
N1_188 <= N0_332;
N1_189 <= N0_333;
N1_190 <= N0_334;
N1_191 <= N0_335;
N1_192 <= N0_336;
N1_193 <= N0_337;
N1_194 <= N0_338;
N1_195 <= N0_339;
N1_196 <= N0_340;
N1_197 <= N0_341;
N1_198 <= N0_342;
N1_199 <= N0_343;
N1_200 <= N0_344;
N1_201 <= N0_345;
N1_202 <= N0_346;
N1_203 <= N0_347;
N1_204 <= N0_348;
N1_205 <= N0_349;
N1_206 <= N0_350;
N1_207 <= N0_351;
N1_208 <= N0_352;
N1_209 <= N0_353;
N1_210 <= N0_354;
N1_211 <= N0_355;
N1_212 <= N0_356;
N1_213 <= N0_357;
N1_214 <= N0_358;
N1_215 <= N0_359;
N2_0 <= N1_0;
N2_1 <= N1_1;
N2_2 <= N1_2;
N2_3 <= N1_3;
N2_4 <= N1_4;
N2_5 <= N1_5;
N2_6 <= N1_6;
N2_7 <= N1_7;
N2_8 <= N1_8;
N2_9 <= N1_9;
N2_10 <= N1_10;
N2_11 <= N1_11;
N2_12 <= N1_12;
N2_13 <= N1_13;
N2_14 <= N1_14;
N2_15 <= N1_15;
N2_16 <= N1_16;
N2_17 <= N1_17;
N2_18 <= N1_18;
N2_19 <= N1_19;
N2_20 <= N1_20;
N2_21 <= N1_21;
N2_22 <= N1_22;
N2_23 <= N1_23;
N2_24 <= N1_24;
N2_25 <= N1_25;
N2_26 <= N1_26;
N2_27 <= N1_27;
N2_28 <= N1_28;
N2_29 <= N1_29;
N2_30 <= N1_30;
N2_31 <= N1_31;
N2_32 <= N1_32;
N2_33 <= N1_33;
N2_34 <= N1_34;
H12 : HA PORT MAP(N1_35,N1_36,H2_0,C2_0);
N2_35 <= N1_37;
N2_36 <= N1_38;
N2_37 <= N1_39;
N2_38 <= N1_40;
N2_39 <= N1_41;
H13 : HA PORT MAP(N1_42,N1_43,H2_1,C2_1);
N2_40 <= N1_44;
N2_41 <= N1_45;
N2_42 <= N1_46;
N2_43 <= N1_47;
F40 : FA PORT MAP(N1_48,N1_49,N1_50,F2_0,C2_2);
H14 : HA PORT MAP(N1_51,N1_52,H2_2,C2_3);
N2_44 <= N1_53;
N2_45 <= N1_54;
N2_46 <= N1_55;
F41 : FA PORT MAP(N1_56,N1_57,N1_58,F2_1,C2_4);
H15 : HA PORT MAP(N1_59,N1_60,H2_3,C2_5);
N2_47 <= N1_61;
N2_48 <= N1_62;
F42 : FA PORT MAP(N1_63,N1_64,N1_65,F2_2,C2_6);
F43 : FA PORT MAP(N1_66,N1_67,N1_68,F2_3,C2_7);
H16 : HA PORT MAP(N1_69,N1_70,H2_4,C2_8);
N2_49 <= N1_71;
F44 : FA PORT MAP(N1_72,N1_73,N1_74,F2_4,C2_9);
F45 : FA PORT MAP(N1_75,N1_76,N1_77,F2_5,C2_10);
H17 : HA PORT MAP(N1_78,N1_79,H2_5,C2_11);
F46 : FA PORT MAP(H1_0,N1_80,N1_81,F2_6,C2_12);
F47 : FA PORT MAP(N1_82,N1_83,N1_84,F2_7,C2_13);
F48 : FA PORT MAP(N1_85,N1_86,N1_87,F2_8,C2_14);
F49 : FA PORT MAP(H1_1,C1_0,N1_88,F2_9,C2_15);
F50 : FA PORT MAP(N1_89,N1_90,N1_91,F2_10,C2_16);
F51 : FA PORT MAP(N1_92,N1_93,N1_94,F2_11,C2_17);
F52 : FA PORT MAP(F1_0,C1_1,H1_2,F2_12,C2_18);
F53 : FA PORT MAP(N1_95,N1_96,N1_97,F2_13,C2_19);
F54 : FA PORT MAP(N1_98,N1_99,N1_100,F2_14,C2_20);
F55 : FA PORT MAP(F1_1,C1_2,H1_3,F2_15,C2_21);
F56 : FA PORT MAP(C1_3,N1_101,N1_102,F2_16,C2_22);
F57 : FA PORT MAP(N1_103,N1_104,N1_105,F2_17,C2_23);
F58 : FA PORT MAP(F1_2,C1_4,F1_3,F2_18,C2_24);
F59 : FA PORT MAP(C1_5,H1_4,N1_106,F2_19,C2_25);
F60 : FA PORT MAP(N1_107,N1_108,N1_109,F2_20,C2_26);
F61 : FA PORT MAP(F1_4,C1_6,F1_5,F2_21,C2_27);
F62 : FA PORT MAP(C1_7,H1_5,C1_8,F2_22,C2_28);
F63 : FA PORT MAP(N1_110,N1_111,N1_112,F2_23,C2_29);
F64 : FA PORT MAP(F1_6,C1_9,F1_7,F2_24,C2_30);
F65 : FA PORT MAP(C1_10,F1_8,C1_11,F2_25,C2_31);
F66 : FA PORT MAP(H1_6,N1_113,N1_114,F2_26,C2_32);
F67 : FA PORT MAP(F1_9,C1_12,F1_10,F2_27,C2_33);
F68 : FA PORT MAP(C1_13,F1_11,C1_14,F2_28,C2_34);
F69 : FA PORT MAP(H1_7,C1_15,N1_115,F2_29,C2_35);
F70 : FA PORT MAP(F1_12,C1_16,F1_13,F2_30,C2_36);
F71 : FA PORT MAP(C1_17,F1_14,C1_18,F2_31,C2_37);
F72 : FA PORT MAP(F1_15,C1_19,N1_116,F2_32,C2_38);
F73 : FA PORT MAP(F1_16,C1_20,F1_17,F2_33,C2_39);
F74 : FA PORT MAP(C1_21,F1_18,C1_22,F2_34,C2_40);
F75 : FA PORT MAP(F1_19,C1_23,N1_117,F2_35,C2_41);
F76 : FA PORT MAP(F1_20,C1_24,F1_21,F2_36,C2_42);
F77 : FA PORT MAP(C1_25,F1_22,C1_26,F2_37,C2_43);
F78 : FA PORT MAP(F1_23,C1_27,N1_118,F2_38,C2_44);
F79 : FA PORT MAP(F1_24,C1_28,F1_25,F2_39,C2_45);
F80 : FA PORT MAP(C1_29,F1_26,C1_30,F2_40,C2_46);
F81 : FA PORT MAP(F1_27,C1_31,N1_119,F2_41,C2_47);
F82 : FA PORT MAP(F1_28,C1_32,F1_29,F2_42,C2_48);
F83 : FA PORT MAP(C1_33,F1_30,C1_34,F2_43,C2_49);
F84 : FA PORT MAP(H1_8,C1_35,N1_120,F2_44,C2_50);
F85 : FA PORT MAP(F1_31,C1_36,F1_32,F2_45,C2_51);
F86 : FA PORT MAP(C1_37,F1_33,C1_38,F2_46,C2_52);
F87 : FA PORT MAP(N1_121,C1_39,N1_122,F2_47,C2_53);
F88 : FA PORT MAP(F1_34,C1_40,F1_35,F2_48,C2_54);
F89 : FA PORT MAP(C1_41,H1_9,C1_42,F2_49,C2_55);
F90 : FA PORT MAP(N1_123,N1_124,N1_125,F2_50,C2_56);
F91 : FA PORT MAP(F1_36,C1_43,F1_37,F2_51,C2_57);
F92 : FA PORT MAP(C1_44,N1_126,C1_45,F2_52,C2_58);
F93 : FA PORT MAP(N1_127,N1_128,N1_129,F2_53,C2_59);
F94 : FA PORT MAP(F1_38,C1_46,H1_10,F2_54,C2_60);
F95 : FA PORT MAP(C1_47,N1_130,N1_131,F2_55,C2_61);
F96 : FA PORT MAP(N1_132,N1_133,N1_134,F2_56,C2_62);
F97 : FA PORT MAP(F1_39,C1_48,N1_135,F2_57,C2_63);
F98 : FA PORT MAP(C1_49,N1_136,N1_137,F2_58,C2_64);
F99 : FA PORT MAP(N1_138,N1_139,N1_140,F2_59,C2_65);
F100 : FA PORT MAP(H1_11,C1_50,N1_141,F2_60,C2_66);
F101 : FA PORT MAP(N1_142,N1_143,N1_144,F2_61,C2_67);
F102 : FA PORT MAP(N1_145,N1_146,N1_147,F2_62,C2_68);
F103 : FA PORT MAP(N1_148,C1_51,N1_149,F2_63,C2_69);
F104 : FA PORT MAP(N1_150,N1_151,N1_152,F2_64,C2_70);
F105 : FA PORT MAP(N1_153,N1_154,N1_155,F2_65,C2_71);
F106 : FA PORT MAP(N1_156,N1_157,N1_158,F2_66,C2_72);
F107 : FA PORT MAP(N1_159,N1_160,N1_161,F2_67,C2_73);
H18 : HA PORT MAP(N1_162,N1_163,H2_6,C2_74);
F108 : FA PORT MAP(N1_164,N1_165,N1_166,F2_68,C2_75);
F109 : FA PORT MAP(N1_167,N1_168,N1_169,F2_69,C2_76);
N2_50 <= N1_170;
F110 : FA PORT MAP(N1_171,N1_172,N1_173,F2_70,C2_77);
H19 : HA PORT MAP(N1_174,N1_175,H2_7,C2_78);
N2_51 <= N1_176;
N2_52 <= N1_177;
F111 : FA PORT MAP(N1_178,N1_179,N1_180,F2_71,C2_79);
N2_53 <= N1_181;
N2_54 <= N1_182;
N2_55 <= N1_183;
H20 : HA PORT MAP(N1_184,N1_185,H2_8,C2_80);
N2_56 <= N1_186;
N2_57 <= N1_187;
N2_58 <= N1_188;
N2_59 <= N1_189;
N2_60 <= N1_190;
N2_61 <= N1_191;
N2_62 <= N1_192;
N2_63 <= N1_193;
N2_64 <= N1_194;
N2_65 <= N1_195;
N2_66 <= N1_196;
N2_67 <= N1_197;
N2_68 <= N1_198;
N2_69 <= N1_199;
N2_70 <= N1_200;
N2_71 <= N1_201;
N2_72 <= N1_202;
N2_73 <= N1_203;
N2_74 <= N1_204;
N2_75 <= N1_205;
N2_76 <= N1_206;
N2_77 <= N1_207;
N2_78 <= N1_208;
N2_79 <= N1_209;
N2_80 <= N1_210;
N2_81 <= N1_211;
N2_82 <= N1_212;
N2_83 <= N1_213;
N2_84 <= N1_214;
N2_85 <= N1_215;
N3_0 <= N2_0;
N3_1 <= N2_1;
N3_2 <= N2_2;
N3_3 <= N2_3;
N3_4 <= N2_4;
N3_5 <= N2_5;
N3_6 <= N2_6;
N3_7 <= N2_7;
N3_8 <= N2_8;
N3_9 <= N2_9;
N3_10 <= N2_10;
N3_11 <= N2_11;
N3_12 <= N2_12;
N3_13 <= N2_13;
N3_14 <= N2_14;
H21 : HA PORT MAP(N2_15,N2_16,H3_0,C3_0);
N3_15 <= N2_17;
N3_16 <= N2_18;
N3_17 <= N2_19;
H22 : HA PORT MAP(N2_20,N2_21,H3_1,C3_1);
N3_18 <= N2_22;
N3_19 <= N2_23;
F112 : FA PORT MAP(N2_24,N2_25,N2_26,F3_0,C3_2);
H23 : HA PORT MAP(N2_27,N2_28,H3_2,C3_3);
N3_20 <= N2_29;
F113 : FA PORT MAP(N2_30,N2_31,N2_32,F3_1,C3_4);
H24 : HA PORT MAP(N2_33,N2_34,H3_3,C3_5);
F114 : FA PORT MAP(H2_0,N2_35,N2_36,F3_2,C3_6);
F115 : FA PORT MAP(N2_37,N2_38,N2_39,F3_3,C3_7);
F116 : FA PORT MAP(H2_1,C2_0,N2_40,F3_4,C3_8);
F117 : FA PORT MAP(N2_41,N2_42,N2_43,F3_5,C3_9);
F118 : FA PORT MAP(F2_0,C2_1,H2_2,F3_6,C3_10);
F119 : FA PORT MAP(N2_44,N2_45,N2_46,F3_7,C3_11);
F120 : FA PORT MAP(F2_1,C2_2,H2_3,F3_8,C3_12);
F121 : FA PORT MAP(C2_3,N2_47,N2_48,F3_9,C3_13);
F122 : FA PORT MAP(F2_2,C2_4,F2_3,F3_10,C3_14);
F123 : FA PORT MAP(C2_5,H2_4,N2_49,F3_11,C3_15);
F124 : FA PORT MAP(F2_4,C2_6,F2_5,F3_12,C3_16);
F125 : FA PORT MAP(C2_7,H2_5,C2_8,F3_13,C3_17);
F126 : FA PORT MAP(F2_6,C2_9,F2_7,F3_14,C3_18);
F127 : FA PORT MAP(C2_10,F2_8,C2_11,F3_15,C3_19);
F128 : FA PORT MAP(F2_9,C2_12,F2_10,F3_16,C3_20);
F129 : FA PORT MAP(C2_13,F2_11,C2_14,F3_17,C3_21);
F130 : FA PORT MAP(F2_12,C2_15,F2_13,F3_18,C3_22);
F131 : FA PORT MAP(C2_16,F2_14,C2_17,F3_19,C3_23);
F132 : FA PORT MAP(F2_15,C2_18,F2_16,F3_20,C3_24);
F133 : FA PORT MAP(C2_19,F2_17,C2_20,F3_21,C3_25);
F134 : FA PORT MAP(F2_18,C2_21,F2_19,F3_22,C3_26);
F135 : FA PORT MAP(C2_22,F2_20,C2_23,F3_23,C3_27);
F136 : FA PORT MAP(F2_21,C2_24,F2_22,F3_24,C3_28);
F137 : FA PORT MAP(C2_25,F2_23,C2_26,F3_25,C3_29);
F138 : FA PORT MAP(F2_24,C2_27,F2_25,F3_26,C3_30);
F139 : FA PORT MAP(C2_28,F2_26,C2_29,F3_27,C3_31);
F140 : FA PORT MAP(F2_27,C2_30,F2_28,F3_28,C3_32);
F141 : FA PORT MAP(C2_31,F2_29,C2_32,F3_29,C3_33);
F142 : FA PORT MAP(F2_30,C2_33,F2_31,F3_30,C3_34);
F143 : FA PORT MAP(C2_34,F2_32,C2_35,F3_31,C3_35);
F144 : FA PORT MAP(F2_33,C2_36,F2_34,F3_32,C3_36);
F145 : FA PORT MAP(C2_37,F2_35,C2_38,F3_33,C3_37);
F146 : FA PORT MAP(F2_36,C2_39,F2_37,F3_34,C3_38);
F147 : FA PORT MAP(C2_40,F2_38,C2_41,F3_35,C3_39);
F148 : FA PORT MAP(F2_39,C2_42,F2_40,F3_36,C3_40);
F149 : FA PORT MAP(C2_43,F2_41,C2_44,F3_37,C3_41);
F150 : FA PORT MAP(F2_42,C2_45,F2_43,F3_38,C3_42);
F151 : FA PORT MAP(C2_46,F2_44,C2_47,F3_39,C3_43);
F152 : FA PORT MAP(F2_45,C2_48,F2_46,F3_40,C3_44);
F153 : FA PORT MAP(C2_49,F2_47,C2_50,F3_41,C3_45);
F154 : FA PORT MAP(F2_48,C2_51,F2_49,F3_42,C3_46);
F155 : FA PORT MAP(C2_52,F2_50,C2_53,F3_43,C3_47);
F156 : FA PORT MAP(F2_51,C2_54,F2_52,F3_44,C3_48);
F157 : FA PORT MAP(C2_55,F2_53,C2_56,F3_45,C3_49);
F158 : FA PORT MAP(F2_54,C2_57,F2_55,F3_46,C3_50);
F159 : FA PORT MAP(C2_58,F2_56,C2_59,F3_47,C3_51);
F160 : FA PORT MAP(F2_57,C2_60,F2_58,F3_48,C3_52);
F161 : FA PORT MAP(C2_61,F2_59,C2_62,F3_49,C3_53);
F162 : FA PORT MAP(F2_60,C2_63,F2_61,F3_50,C3_54);
F163 : FA PORT MAP(C2_64,F2_62,C2_65,F3_51,C3_55);
F164 : FA PORT MAP(F2_63,C2_66,F2_64,F3_52,C3_56);
F165 : FA PORT MAP(C2_67,F2_65,C2_68,F3_53,C3_57);
F166 : FA PORT MAP(F2_66,C2_69,F2_67,F3_54,C3_58);
F167 : FA PORT MAP(C2_70,H2_6,C2_71,F3_55,C3_59);
F168 : FA PORT MAP(F2_68,C2_72,F2_69,F3_56,C3_60);
F169 : FA PORT MAP(C2_73,N2_50,C2_74,F3_57,C3_61);
F170 : FA PORT MAP(F2_70,C2_75,H2_7,F3_58,C3_62);
F171 : FA PORT MAP(C2_76,N2_51,N2_52,F3_59,C3_63);
F172 : FA PORT MAP(F2_71,C2_77,N2_53,F3_60,C3_64);
F173 : FA PORT MAP(C2_78,N2_54,N2_55,F3_61,C3_65);
F174 : FA PORT MAP(H2_8,C2_79,N2_56,F3_62,C3_66);
F175 : FA PORT MAP(N2_57,N2_58,N2_59,F3_63,C3_67);
F176 : FA PORT MAP(N2_60,C2_80,N2_61,F3_64,C3_68);
F177 : FA PORT MAP(N2_62,N2_63,N2_64,F3_65,C3_69);
F178 : FA PORT MAP(N2_65,N2_66,N2_67,F3_66,C3_70);
H25 : HA PORT MAP(N2_68,N2_69,H3_4,C3_71);
F179 : FA PORT MAP(N2_70,N2_71,N2_72,F3_67,C3_72);
N3_21 <= N2_73;
H26 : HA PORT MAP(N2_74,N2_75,H3_5,C3_73);
N3_22 <= N2_76;
N3_23 <= N2_77;
N3_24 <= N2_78;
N3_25 <= N2_79;
N3_26 <= N2_80;
N3_27 <= N2_81;
N3_28 <= N2_82;
N3_29 <= N2_83;
N3_30 <= N2_84;
N3_31 <= N2_85;
N4_0 <= N3_0;
N4_1 <= N3_1;
N4_2 <= N3_2;
N4_3 <= N3_3;
N4_4 <= N3_4;
N4_5 <= N3_5;
N4_6 <= N3_6;
N4_7 <= N3_7;
H27 : HA PORT MAP(N3_8,N3_9,H4_0,C4_0);
N4_8 <= N3_10;
N4_9 <= N3_11;
H28 : HA PORT MAP(N3_12,N3_13,H4_1,C4_1);
N4_10 <= N3_14;
F180 : FA PORT MAP(H3_0,N3_15,N3_16,F4_0,C4_2);
N4_11 <= N3_17;
F181 : FA PORT MAP(H3_1,C3_0,N3_18,F4_1,C4_3);
N4_12 <= N3_19;
F182 : FA PORT MAP(F3_0,C3_1,H3_2,F4_2,C4_4);
N4_13 <= N3_20;
F183 : FA PORT MAP(F3_1,C3_2,H3_3,F4_3,C4_5);
N4_14 <= C3_3;
F184 : FA PORT MAP(F3_2,C3_4,F3_3,F4_4,C4_6);
N4_15 <= C3_5;
F185 : FA PORT MAP(F3_4,C3_6,F3_5,F4_5,C4_7);
N4_16 <= C3_7;
F186 : FA PORT MAP(F3_6,C3_8,F3_7,F4_6,C4_8);
N4_17 <= C3_9;
F187 : FA PORT MAP(F3_8,C3_10,F3_9,F4_7,C4_9);
N4_18 <= C3_11;
F188 : FA PORT MAP(F3_10,C3_12,F3_11,F4_8,C4_10);
N4_19 <= C3_13;
F189 : FA PORT MAP(F3_12,C3_14,F3_13,F4_9,C4_11);
N4_20 <= C3_15;
F190 : FA PORT MAP(F3_14,C3_16,F3_15,F4_10,C4_12);
N4_21 <= C3_17;
F191 : FA PORT MAP(F3_16,C3_18,F3_17,F4_11,C4_13);
N4_22 <= C3_19;
F192 : FA PORT MAP(F3_18,C3_20,F3_19,F4_12,C4_14);
N4_23 <= C3_21;
F193 : FA PORT MAP(F3_20,C3_22,F3_21,F4_13,C4_15);
N4_24 <= C3_23;
F194 : FA PORT MAP(F3_22,C3_24,F3_23,F4_14,C4_16);
N4_25 <= C3_25;
F195 : FA PORT MAP(F3_24,C3_26,F3_25,F4_15,C4_17);
N4_26 <= C3_27;
F196 : FA PORT MAP(F3_26,C3_28,F3_27,F4_16,C4_18);
N4_27 <= C3_29;
F197 : FA PORT MAP(F3_28,C3_30,F3_29,F4_17,C4_19);
N4_28 <= C3_31;
F198 : FA PORT MAP(F3_30,C3_32,F3_31,F4_18,C4_20);
N4_29 <= C3_33;
F199 : FA PORT MAP(F3_32,C3_34,F3_33,F4_19,C4_21);
N4_30 <= C3_35;
F200 : FA PORT MAP(F3_34,C3_36,F3_35,F4_20,C4_22);
N4_31 <= C3_37;
F201 : FA PORT MAP(F3_36,C3_38,F3_37,F4_21,C4_23);
N4_32 <= C3_39;
F202 : FA PORT MAP(F3_38,C3_40,F3_39,F4_22,C4_24);
N4_33 <= C3_41;
F203 : FA PORT MAP(F3_40,C3_42,F3_41,F4_23,C4_25);
N4_34 <= C3_43;
F204 : FA PORT MAP(F3_42,C3_44,F3_43,F4_24,C4_26);
N4_35 <= C3_45;
F205 : FA PORT MAP(F3_44,C3_46,F3_45,F4_25,C4_27);
N4_36 <= C3_47;
F206 : FA PORT MAP(F3_46,C3_48,F3_47,F4_26,C4_28);
N4_37 <= C3_49;
F207 : FA PORT MAP(F3_48,C3_50,F3_49,F4_27,C4_29);
N4_38 <= C3_51;
F208 : FA PORT MAP(F3_50,C3_52,F3_51,F4_28,C4_30);
N4_39 <= C3_53;
F209 : FA PORT MAP(F3_52,C3_54,F3_53,F4_29,C4_31);
N4_40 <= C3_55;
F210 : FA PORT MAP(F3_54,C3_56,F3_55,F4_30,C4_32);
N4_41 <= C3_57;
F211 : FA PORT MAP(F3_56,C3_58,F3_57,F4_31,C4_33);
N4_42 <= C3_59;
F212 : FA PORT MAP(F3_58,C3_60,F3_59,F4_32,C4_34);
N4_43 <= C3_61;
F213 : FA PORT MAP(F3_60,C3_62,F3_61,F4_33,C4_35);
N4_44 <= C3_63;
F214 : FA PORT MAP(F3_62,C3_64,F3_63,F4_34,C4_36);
N4_45 <= C3_65;
F215 : FA PORT MAP(F3_64,C3_66,F3_65,F4_35,C4_37);
N4_46 <= C3_67;
F216 : FA PORT MAP(F3_66,C3_68,H3_4,F4_36,C4_38);
N4_47 <= C3_69;
F217 : FA PORT MAP(F3_67,C3_70,N3_21,F4_37,C4_39);
N4_48 <= C3_71;
F218 : FA PORT MAP(H3_5,C3_72,N3_22,F4_38,C4_40);
N4_49 <= N3_23;
F219 : FA PORT MAP(N3_24,C3_73,N3_25,F4_39,C4_41);
N4_50 <= N3_26;
H29 : HA PORT MAP(N3_27,N3_28,H4_2,C4_42);
N4_51 <= N3_29;
N4_52 <= N3_30;
N4_53 <= N3_31;
N5_0 <= N4_0;
N5_1 <= N4_1;
N5_2 <= N4_2;
H30 : HA PORT MAP(N4_3,N4_4,H5_0,C5_0);
N5_3 <= N4_5;
H31 : HA PORT MAP(N4_6,N4_7,H5_1,C5_1);
F220 : FA PORT MAP(H4_0,N4_8,N4_9,F5_0,C5_2);
F221 : FA PORT MAP(H4_1,C4_0,N4_10,F5_1,C5_3);
F222 : FA PORT MAP(F4_0,C4_1,N4_11,F5_2,C5_4);
F223 : FA PORT MAP(F4_1,C4_2,N4_12,F5_3,C5_5);
F224 : FA PORT MAP(F4_2,C4_3,N4_13,F5_4,C5_6);
F225 : FA PORT MAP(F4_3,C4_4,N4_14,F5_5,C5_7);
F226 : FA PORT MAP(F4_4,C4_5,N4_15,F5_6,C5_8);
F227 : FA PORT MAP(F4_5,C4_6,N4_16,F5_7,C5_9);
F228 : FA PORT MAP(F4_6,C4_7,N4_17,F5_8,C5_10);
F229 : FA PORT MAP(F4_7,C4_8,N4_18,F5_9,C5_11);
F230 : FA PORT MAP(F4_8,C4_9,N4_19,F5_10,C5_12);
F231 : FA PORT MAP(F4_9,C4_10,N4_20,F5_11,C5_13);
F232 : FA PORT MAP(F4_10,C4_11,N4_21,F5_12,C5_14);
F233 : FA PORT MAP(F4_11,C4_12,N4_22,F5_13,C5_15);
F234 : FA PORT MAP(F4_12,C4_13,N4_23,F5_14,C5_16);
F235 : FA PORT MAP(F4_13,C4_14,N4_24,F5_15,C5_17);
F236 : FA PORT MAP(F4_14,C4_15,N4_25,F5_16,C5_18);
F237 : FA PORT MAP(F4_15,C4_16,N4_26,F5_17,C5_19);
F238 : FA PORT MAP(F4_16,C4_17,N4_27,F5_18,C5_20);
F239 : FA PORT MAP(F4_17,C4_18,N4_28,F5_19,C5_21);
F240 : FA PORT MAP(F4_18,C4_19,N4_29,F5_20,C5_22);
F241 : FA PORT MAP(F4_19,C4_20,N4_30,F5_21,C5_23);
F242 : FA PORT MAP(F4_20,C4_21,N4_31,F5_22,C5_24);
F243 : FA PORT MAP(F4_21,C4_22,N4_32,F5_23,C5_25);
F244 : FA PORT MAP(F4_22,C4_23,N4_33,F5_24,C5_26);
F245 : FA PORT MAP(F4_23,C4_24,N4_34,F5_25,C5_27);
F246 : FA PORT MAP(F4_24,C4_25,N4_35,F5_26,C5_28);
F247 : FA PORT MAP(F4_25,C4_26,N4_36,F5_27,C5_29);
F248 : FA PORT MAP(F4_26,C4_27,N4_37,F5_28,C5_30);
F249 : FA PORT MAP(F4_27,C4_28,N4_38,F5_29,C5_31);
F250 : FA PORT MAP(F4_28,C4_29,N4_39,F5_30,C5_32);
F251 : FA PORT MAP(F4_29,C4_30,N4_40,F5_31,C5_33);
F252 : FA PORT MAP(F4_30,C4_31,N4_41,F5_32,C5_34);
F253 : FA PORT MAP(F4_31,C4_32,N4_42,F5_33,C5_35);
F254 : FA PORT MAP(F4_32,C4_33,N4_43,F5_34,C5_36);
F255 : FA PORT MAP(F4_33,C4_34,N4_44,F5_35,C5_37);
F256 : FA PORT MAP(F4_34,C4_35,N4_45,F5_36,C5_38);
F257 : FA PORT MAP(F4_35,C4_36,N4_46,F5_37,C5_39);
F258 : FA PORT MAP(F4_36,C4_37,N4_47,F5_38,C5_40);
F259 : FA PORT MAP(F4_37,C4_38,N4_48,F5_39,C5_41);
F260 : FA PORT MAP(F4_38,C4_39,N4_49,F5_40,C5_42);
F261 : FA PORT MAP(F4_39,C4_40,N4_50,F5_41,C5_43);
F262 : FA PORT MAP(H4_2,C4_41,N4_51,F5_42,C5_44);
F263 : FA PORT MAP(N4_52,C4_42,N4_53,F5_43,open);
H32 : HA PORT MAP(N5_0,N5_1,Y(0),Co_0);
H33 : HA PORT MAP(N5_2,Co_0,Y(1),Co_1);
F264 : FA PORT MAP(H5_0,N5_3,Co_1,Y(2),Co_2);
F265 : FA PORT MAP(H5_1,C5_0,Co_2,Y(3),Co_3);
F266 : FA PORT MAP(F5_0,C5_1,Co_3,Y(4),Co_4);
F267 : FA PORT MAP(F5_1,C5_2,Co_4,Y(5),Co_5);
F268 : FA PORT MAP(F5_2,C5_3,Co_5,Y(6),Co_6);
F269 : FA PORT MAP(F5_3,C5_4,Co_6,Y(7),Co_7);
F270 : FA PORT MAP(F5_4,C5_5,Co_7,Y(8),Co_8);
F271 : FA PORT MAP(F5_5,C5_6,Co_8,Y(9),Co_9);
F272 : FA PORT MAP(F5_6,C5_7,Co_9,Y(10),Co_10);
F273 : FA PORT MAP(F5_7,C5_8,Co_10,Y(11),Co_11);
F274 : FA PORT MAP(F5_8,C5_9,Co_11,Y(12),Co_12);
F275 : FA PORT MAP(F5_9,C5_10,Co_12,Y(13),Co_13);
F276 : FA PORT MAP(F5_10,C5_11,Co_13,Y(14),Co_14);
F277 : FA PORT MAP(F5_11,C5_12,Co_14,Y(15),Co_15);
F278 : FA PORT MAP(F5_12,C5_13,Co_15,Y(16),Co_16);
F279 : FA PORT MAP(F5_13,C5_14,Co_16,Y(17),Co_17);
F280 : FA PORT MAP(F5_14,C5_15,Co_17,Y(18),Co_18);
F281 : FA PORT MAP(F5_15,C5_16,Co_18,Y(19),Co_19);
F282 : FA PORT MAP(F5_16,C5_17,Co_19,Y(20),Co_20);
F283 : FA PORT MAP(F5_17,C5_18,Co_20,Y(21),Co_21);
F284 : FA PORT MAP(F5_18,C5_19,Co_21,Y(22),Co_22);
F285 : FA PORT MAP(F5_19,C5_20,Co_22,Y(23),Co_23);
F286 : FA PORT MAP(F5_20,C5_21,Co_23,Y(24),Co_24);
F287 : FA PORT MAP(F5_21,C5_22,Co_24,Y(25),Co_25);
F288 : FA PORT MAP(F5_22,C5_23,Co_25,Y(26),Co_26);
F289 : FA PORT MAP(F5_23,C5_24,Co_26,Y(27),Co_27);
F290 : FA PORT MAP(F5_24,C5_25,Co_27,Y(28),Co_28);
F291 : FA PORT MAP(F5_25,C5_26,Co_28,Y(29),Co_29);
F292 : FA PORT MAP(F5_26,C5_27,Co_29,Y(30),Co_30);
F293 : FA PORT MAP(F5_27,C5_28,Co_30,Y(31),Co_31);
F294 : FA PORT MAP(F5_28,C5_29,Co_31,Y(32),Co_32);
F295 : FA PORT MAP(F5_29,C5_30,Co_32,Y(33),Co_33);
F296 : FA PORT MAP(F5_30,C5_31,Co_33,Y(34),Co_34);
F297 : FA PORT MAP(F5_31,C5_32,Co_34,Y(35),Co_35);
F298 : FA PORT MAP(F5_32,C5_33,Co_35,Y(36),Co_36);
F299 : FA PORT MAP(F5_33,C5_34,Co_36,Y(37),Co_37);
F300 : FA PORT MAP(F5_34,C5_35,Co_37,Y(38),Co_38);
F301 : FA PORT MAP(F5_35,C5_36,Co_38,Y(39),Co_39);
F302 : FA PORT MAP(F5_36,C5_37,Co_39,Y(40),Co_40);
F303 : FA PORT MAP(F5_37,C5_38,Co_40,Y(41),Co_41);
F304 : FA PORT MAP(F5_38,C5_39,Co_41,Y(42),Co_42);
F305 : FA PORT MAP(F5_39,C5_40,Co_42,Y(43),Co_43);
F306 : FA PORT MAP(F5_40,C5_41,Co_43,Y(44),Co_44);
F307 : FA PORT MAP(F5_41,C5_42,Co_44,Y(45),Co_45);
F308 : FA PORT MAP(F5_42,C5_43,Co_45,Y(46),Co_46);
F309 : FA PORT MAP(F5_43,C5_44,Co_46,Y(47),open);
END behavior;